** sch_path: /foss/designs/SAR_ADC_IHP/xschem/dac_icms_cell/testbenches/tb_capacitor.sch
**.subckt tb_capacitor
V7 sample GND PULSE( 0 1.8 0 10p 10p 5n 10n 1)
x10 VDD sample net1 GND inverter_lv W_P=1.0u L_P=0.13u W_N=1.0u L_N=0.13u n=16
V2 vin GND 1.7
V3 vcm GND 0.9
V4 VDD GND 1.8
C1 vcbot vctop 20f m=64
V1 vcbot net4 0
V5 vcbot net5 0
V6 sample_n net1 0
V8 sample net11 0
XM1 vin sample_s net3 GND sg13_lv_nmos w=0.15u l=0.13u ng=1 m=64
XM2 vin sample_n net2 VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=64
XM3 net3 sample_n net3 GND sg13_lv_nmos w=0.15u l=0.13u ng=1 m=32
XM4 net2 sample_s net2 VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=32
x1 VDD net1 sample_s GND inverter_lv W_P=1.0u L_P=0.13u W_N=1.0u L_N=0.13u n=16
V9 net10 vcm 0
XM5 net2 GND net4 VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=32
XM6 net3 VDD net5 GND sg13_lv_nmos w=0.15u l=0.13u ng=1 m=32
V10 vctop net8 0
V11 vctop net9 0
XM7 vcm sample_s net7 GND sg13_lv_nmos w=0.15u l=0.13u ng=1 m=64
XM8 vcm sample_n net6 VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=64
XM9 net7 sample_n net7 GND sg13_lv_nmos w=0.15u l=0.13u ng=1 m=32
XM10 net6 sample_s net6 VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=32
XM11 net6 GND net8 VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=32
XM12 net7 VDD net9 GND sg13_lv_nmos w=0.15u l=0.13u ng=1 m=32
**** begin user architecture code


.param temp=27
.param W_P = 1.0u
.param L_P = 0.13u
.param W_N = 1.0u
.param L_N = 0.13u
.options savecurrents klu method=gear reltol=1e-2 abstol=1e-15 gmin=1e-10
.control

* Transient Analysis
tran 100p 20n

*plot {d0} {d1 + 4} {d2 + 8} {d3 + 12} {d4 + 16} {d5 + 20} {d6 + 24} {d7 + 28} {d8 + 32} {d9 + 36} {d10 + 40} {d11 + 44}
*plot {b0} {b1 + 4} {b2 + 8} {b3 + 12} {b4 + 16} {b5 + 20} {b6 + 24} {b7 + 28} {b8 + 32} {b9 + 36} {b10 + 40} {b11 + 44}
*plot {clk} {comp_in + 2} {sample + 4}
plot vctop vcbot sample
plot {vctop-vcbot} sample
plot i(v1) i(v5)
*plot x3.x14.net1-vctop x3.x18.vcap-vcbot

.endc




** IHP models
.lib cornerMOSlv.lib mos_tt
.lib cornerMOShv.lib mos_tt
.lib cornerHBT.lib hbt_typ
.lib cornerRES.lib res_typ
.include /foss/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice


**** end user architecture code
**.ends

* expanding   symbol:  inverter/inverter_lv.sym # of pins=4
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/inverter/inverter_lv.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/inverter/inverter_lv.sch
.subckt inverter_lv VDD vin vout VSS  W_P=3.0u L_P=0.13u W_N=1.0u L_N=0.13u n=1
*.ipin vin
*.iopin VDD
*.iopin VSS
*.opin vout
XM1 vout vin VDD VDD sg13_lv_pmos w=W_P l=L_P ng=1 m=n
XM2 vout vin VSS VSS sg13_lv_nmos w=W_N l=L_N ng=1 m=n
.ends

.GLOBAL GND
.end
