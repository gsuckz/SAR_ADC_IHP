** sch_path: /foss/designs/SAR_ADC_IHP/xschem/comparator/pulse_gen/testbench/tb_pgen.sch
**.subckt tb_pgen
x1 VDD GND GND comp PULSEN VTUNE pgen
VDD VDD GND 1.5
VDD1 VTUNE GND 1.1
VDD2 comp GND PULSE(0 1.5 50n 10p 10p 10n 100n)
x6 PULSEN VDD VSS PULSE sg13g2_inv_2
VDD3 VSS GND 0
**** begin user architecture code

.lib cornerMOSlv.lib mos_tt
.lib cornerMOShv.lib mos_tt
.lib cornerRES.lib res_typ
.include /foss/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice



.param temp=27
*.options savecurrents reltol=1e-3 abstol=1e-12 gmin=1e-15
.control
save all

tran 40p 450n

* Plotting
plot v(comp) {v(x1.vx) + 2} {v(PULSE)  +4} {x1.READY + 6} {v(PULSEN) + 8}

.endc

**** end user architecture code
**.ends

* expanding   symbol:  comparator/pulse_gen/pgen.sym # of pins=6
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/comparator/pulse_gen/pgen.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/comparator/pulse_gen/pgen.sch
.subckt pgen VDD in2 VSS in1 PULSE_n VTUNE
*.iopin VDD
*.iopin in2
*.iopin in1
*.iopin VSS
*.iopin VTUNE
*.iopin PULSE_n
XM1 READY in1 VSS VSS sg13_lv_nmos w=2u l=0.13u ng=1 m=1
XM2 READY vx_n VDD VDD sg13_lv_pmos w=2u l=0.13u ng=1 m=1
XM4 vx PULSE_n net4 VDD sg13_lv_pmos w=2u l=0.13u ng=1 m=1
x46 vxs READY VDD VSS PULSE_n sg13g2_or2_2
x6 vxs VDD VSS vx_n sg13g2_inv_2
XM3 READY in2 VSS VSS sg13_lv_nmos w=2u l=0.13u ng=1 m=1
XM5 vx READY VSS VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM7 net4 VTUNE VDD VDD sg13_lv_pmos w=2u l=0.13u ng=1 m=1
XM6 net3 vx VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM8 net2 vx net1 VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM9 net2 vx net3 VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM10 net1 vx VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM11 VDD net2 net1 VDD sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM12 VSS net2 net3 VSS sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
x1 net2 VDD VSS vxs sg13g2_inv_2
.ends

.GLOBAL GND
.GLOBAL VDD
.GLOBAL VTUNE
.GLOBAL comp
.end
