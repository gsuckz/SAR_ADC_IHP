** sch_path: /foss/pdks/ihp-sg13g2/libs.tech/xschem/sg13g2_tests/tran_mim_cap.sch
**.subckt tran_mim_cap
I1 0 G pwl 0 0 1000n 0 1010n 100n
R1 G REF 1G m=1
I3 0 G2 pwl 0 0 1000n 0 1010n 100n
R3 G2 REF 1G m=1
C1 G2 0 0.07452p m=1
V1 REF 0 -2
XC2 G 0 cap_cmim w=7.0e-6 l=7.0e-6 m=1
**** begin user architecture code


.control
save all
tran 10n 6u
write test_mim_cap.raw
.endc



.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerCAP.lib cap_typ

**** end user architecture code
**.ends
.end
