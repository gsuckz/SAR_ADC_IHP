** sch_path: /foss/designs/SAR_ADC_IHP/xschem/untitled-1.sch
**.subckt untitled-1
I0 GND v1 PULSE(0 1m 0 10p 10p 1n 4n)
R1 v1 GND 1k m=1
I1 v1 GND PULSE(0 1m 2n 10p 10p 1n 4n)
**** begin user architecture code


.param temp=27
*.options savecurrents reltol=1e-3 abstol=1e-12 gmin=1e-15
.control
save all

tran 1p 40n

* Plotting
plot v1

.endc

**** end user architecture code
**.ends
.GLOBAL GND
.end
