** sch_path: /foss/designs/SAR_ADC_IHP/xschem/dac_icms_cell/testbenches/tb_unit_cell_logic_reg_tran.sch
**.subckt tb_unit_cell_logic_reg_tran
x1 bit net1 GND d vdd top unit_cell W_P_SPDT=1.0u L_P_SPDT=0.13u W_N_SPDT=1.0u L_N_SPDT=0.13u Cu=20f n=32
V1 vdd GND 1.8
V2 clk GND PULSE( 0 1.8 0 10p 10p 2n 4n)
V3 vcm GND 0.9
V4 comp_in GND 0
S1 top vcm s GND SW1
V5 s GND PULSE(-10 10 0 10p 10p 10n 20n 1)
S2 net2 net1 s GND SW1
S3 vcm net1 GND s SW1
V6 net2 GND 1
x18 clk p_dec vdd comp_in vdd bit GND d bit_cell
V7 p_dec GND PULSE(1.8 0 0 10p 10p 15n 20n 1)
x2 bit net3 GND d vdd top_n unit_cell_n W_P_SPDT=1.0u L_P_SPDT=0.13u W_N_SPDT=1.0u L_N_SPDT=0.13u Cu=20f n=32
S4 top_n vcm s GND SW1
S5 GND net3 s GND SW1
S6 vcm net3 GND s SW1
x3 clk d vdd comp_in vdd bit2 GND d2 bit_cell
x4 bit2 net4 GND d2 vdd top unit_cell W_P_SPDT=1.0u L_P_SPDT=0.13u W_N_SPDT=1.0u L_N_SPDT=0.13u Cu=20f n=16
S7 top vcm s GND SW1
S8 net5 net4 s GND SW1
S9 vcm net4 GND s SW1
V8 net5 GND 1
x5 bit2 net6 GND d2 vdd top_n unit_cell_n W_P_SPDT=1.0u L_P_SPDT=0.13u W_N_SPDT=1.0u L_N_SPDT=0.13u Cu=20f n=16
S10 top_n vcm s GND SW1
S11 GND net6 s GND SW1
S12 vcm net6 GND s SW1
x6 bit3 net7 GND d3 vdd top2 unit_cell W_P_SPDT=1.0u L_P_SPDT=0.13u W_N_SPDT=1.0u L_N_SPDT=0.13u Cu=20f n=32
S13 top2 vcm s GND SW1
S14 net8 net7 s GND SW1
S15 vcm net7 GND s SW1
V9 net8 GND 1
x7 bit3 net9 GND d3 vdd top_n2 unit_cell_n W_P_SPDT=1.0u L_P_SPDT=0.13u W_N_SPDT=1.0u L_N_SPDT=0.13u Cu=20f n=32
S16 top_n2 vcm s GND SW1
S17 GND net9 s GND SW1
S18 vcm net9 GND s SW1
x8 bit4 net10 GND d4 vdd top2 unit_cell W_P_SPDT=1.0u L_P_SPDT=0.13u W_N_SPDT=1.0u L_N_SPDT=0.13u Cu=20f n=16
S19 top2 vcm s GND SW1
S20 net11 net10 s GND SW1
S21 vcm net10 GND s SW1
V10 net11 GND 1
x9 bit4 net12 GND d4 vdd top_n2 unit_cell_n W_P_SPDT=1.0u L_P_SPDT=0.13u W_N_SPDT=1.0u L_N_SPDT=0.13u Cu=20f n=16
S22 top_n2 vcm s GND SW1
S23 GND net12 s GND SW1
S24 vcm net12 GND s SW1
C1 top2 top 20f m=22
C2 top_n2 top_n 20f m=22
x10 clk d2 vdd comp_in vdd bit3 GND d3 bit_cell
x11 clk d3 vdd comp_in vdd bit4 GND d4 bit_cell
C3 top2 net7 20f m=16
C4 top_n2 net9 20f m=16
**** begin user architecture code


.param temp=27
.param W_P = 1.0u
.param L_P = 0.13u
.param W_N = 1.0u
.param L_N = 0.13u
*.options savecurrents klu method=gear reltol=1e-2 abstol=1e-15 gmin=1e-15
.control

* Transient Analysis
tran 10p 40n

plot top {bit +2} {d +4} {s + 6}
plot i(V2) i(V3) i(V6)
plot clk comp_in+3 p_dec+6
plot top top_n

.endc




** IHP models
.lib cornerMOSlv.lib mos_tt
.lib cornerMOShv.lib mos_tt
.lib cornerHBT.lib hbt_typ
.lib cornerRES.lib res_typ
.include /foss/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice


**** end user architecture code
**.ends

* expanding   symbol:  dac_icms_cell/unit_cell.sym # of pins=6
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/dac_icms_cell/unit_cell.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/dac_icms_cell/unit_cell.sch
.subckt unit_cell B A VSS D VDD vtop  W_P_SPDT=1.0u L_P_SPDT=0.13u W_N_SPDT=1.0u L_N_SPDT=0.13u Cu=8f n=1
*.iopin VSS
*.iopin A
*.iopin VDD
*.ipin D
*.iopin B
*.iopin vtop
x1 VDD D VSS vcap B A dac_switch W_P_TG=3.0u L_P_TG=0.13u W_N_TG=1.0u L_N_TG=0.13u n=n
C1 vcap vtop Cu m=n
.ends


* expanding   symbol:  logic/bit_cell.sym # of pins=8
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/logic/bit_cell.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/logic/bit_cell.sch
.subckt bit_cell clk p_bit_dec reset comp_in VDD bit VSS dec
*.iopin p_bit_dec
*.iopin clk
*.iopin reset
*.iopin comp_in
*.iopin VDD
*.iopin VSS
*.iopin bit
*.iopin dec
x1 VDD net2 net4 VSS net5 net1 SR_latch W_P_SR=1.0u L_P_SR=0.13u W_N_SR=1.0u L_N_SR=0.13u
x23 net6 n_dec VDD VSS net1 sg13g2_and2_1
x14 n_dec comp_in VDD VSS net2 sg13g2_and2_1
x30 comp_in VDD VSS net6 sg13g2_inv_2
x53 clk p_bit_dec net3 n_dec reset VDD VSS sg13g2_dfrbp_1
* noconn #net4
x2 VDD net5 net7 VSS buffer_lv W_P_INV=3.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x3 VDD net3 net8 VSS buffer_lv W_P_INV=3.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x4 VDD net8 dec VSS buffer_lv W_P_INV=10.0u L_P_INV=0.13u W_N_INV=10.0u L_N_INV=0.13u
x5 VDD net7 bit VSS buffer_lv W_P_INV=10.0u L_P_INV=0.13u W_N_INV=10.0u L_N_INV=0.13u
.ends


* expanding   symbol:  dac_icms_cell/unit_cell_n.sym # of pins=6
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/dac_icms_cell/unit_cell_n.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/dac_icms_cell/unit_cell_n.sch
.subckt unit_cell_n B A VSS D VDD vtop  W_P_SPDT=1.0u L_P_SPDT=0.13u W_N_SPDT=1.0u L_N_SPDT=0.13u Cu=8f n=1
*.iopin VSS
*.iopin A
*.iopin VDD
*.ipin D
*.iopin B
*.iopin vtop
x1 VDD D VSS net1 B A dac_switch_n W_P_TG=3.0u L_P_TG=0.13u W_N_TG=1.0u L_N_TG=0.13u n=n
C1 net1 vtop cu m=n
.ends


* expanding   symbol:  dac_icms_cell/dac_switch.sym # of pins=6
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/dac_icms_cell/dac_switch.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/dac_icms_cell/dac_switch.sch
.subckt dac_switch VDD di_spdt_ctrl VSS v_c v_b v_a  W_P_TG=3.0u L_P_TG=0.13u W_N_TG=1.0u L_N_TG=0.13u n=1
*.iopin v_a
*.iopin v_c
*.iopin VDD
*.iopin VSS
*.ipin di_spdt_ctrl
*.iopin v_b
x1 VDD di_spdt_ctrl_n VSS net2 v_a di_spdt_ctrl transmission_gate_lv_w_dummy W_P=W_P_TG L_P=L_P_TG W_N=W_N_TG L_N=L_N_TG
+ W_P_D=1.0u L_P_D=0.13u W_N_D=1.0u L_N_D=0.13u n=n
x8 VDD di_spdt_ctrl di_spdt_ctrl_n VSS inverter_lv W_P=W_P_TG L_P=L_P_TG W_N=W_N_TG L_N=L_N_TG n=n
XM1 net1 v_b VSS VSS sg13_lv_nmos w=0.5u l=0.2u ng=1 m=n
XM3 net1 v_b VDD VDD sg13_lv_pmos w=1u l=0.2u ng=1 m=n
x2 VDD di_spdt_ctrl VSS net3 net1 di_spdt_ctrl_n transmission_gate_lv_w_dummy W_P=W_P_TG L_P=L_P_TG W_N=W_N_TG L_N=L_N_TG
+ W_P_D=1.0u L_P_D=0.13u W_N_D=1.0u L_N_D=0.13u n=n
V1 v_c net2 0
V2 v_c net3 0
.ends


* expanding   symbol:  comparator/SR_latch/SR_latch.sym # of pins=6
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/comparator/SR_latch/SR_latch.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/comparator/SR_latch/SR_latch.sch
.subckt SR_latch VDD S Qn VSS Q R  W_P_SR=1.0u L_P_SR=0.13u W_N_SR=1.0u L_N_SR=0.13u
*.iopin VDD
*.opin Q
*.iopin VSS
*.ipin S
*.ipin R
*.opin Qn
x1 VDD Q R Qn VSS NOR_gate W_P=W_P_SR L_P=L_P_SR W_N=W_N_SR L_N=L_N_SR
x2 VDD Qn Q S VSS NOR_gate W_P=W_P_SR L_P=L_P_SR W_N=W_N_SR L_N=L_N_SR
.ends


* expanding   symbol:  buffer/buffer_lv.sym # of pins=4
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/buffer/buffer_lv.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/buffer/buffer_lv.sch
.subckt buffer_lv VDD vin vout VSS  W_P_INV=3.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
*.ipin vin
*.iopin VDD
*.iopin VSS
*.opin vout
x1 VDD vin net1 VSS inverter_lv W_P=W_P_INV L_P=L_P_INV W_N=W_N_INV L_N=L_N_INV n=1
x2 VDD net1 vout VSS inverter_lv W_P=W_P_INV L_P=L_P_INV W_N=W_N_INV L_N=L_N_INV n=1
.ends


* expanding   symbol:  dac_icms_cell/dac_switch_n.sym # of pins=6
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/dac_icms_cell/dac_switch_n.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/dac_icms_cell/dac_switch_n.sch
.subckt dac_switch_n VDD di_spdt_ctrl VSS v_c v_b v_a  W_P_TG=3.0u L_P_TG=0.13u W_N_TG=1.0u L_N_TG=0.13u n=1
*.iopin v_a
*.iopin v_c
*.iopin VDD
*.iopin VSS
*.ipin di_spdt_ctrl
*.iopin v_b
x1 VDD di_spdt_ctrl_n VSS v_c v_a di_spdt_ctrl transmission_gate_lv_wo_dummy W_P=W_P_TG L_P=L_P_TG W_N=W_N_TG L_N=L_N_TG
x8 VDD di_spdt_ctrl di_spdt_ctrl_n VSS inverter_lv W_P=W_P_TG L_P=L_P_TG W_N=W_N_TG L_N=L_N_TG n=n
XM1 net1 net2 VSS VSS sg13_lv_nmos w=0.5u l=0.2u ng=1 m=n
XM3 net1 net2 VDD VDD sg13_lv_pmos w=1u l=0.2u ng=1 m=n
x2 VDD di_spdt_ctrl VSS v_c net1 di_spdt_ctrl_n transmission_gate_lv_w_dummy W_P=W_P_TG L_P=L_P_TG W_N=W_N_TG L_N=L_N_TG
+ W_P_D=1.0u L_P_D=0.13u W_N_D=1.0u L_N_D=0.13u n=n
XM2 net2 v_b VSS VSS sg13_lv_nmos w=0.5u l=0.2u ng=1 m=10
XM4 net2 v_b VDD VDD sg13_lv_pmos w=1u l=0.2u ng=1 m=10
.ends


* expanding   symbol:  transmission_gate/transmission_gate_lv_w_dummy.sym # of pins=6
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/transmission_gate/transmission_gate_lv_w_dummy.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/transmission_gate/transmission_gate_lv_w_dummy.sch
.subckt transmission_gate_lv_w_dummy VDD di_tg_ctrl VSS v_b v_a di_tg_ctrl_n  W_P=2.0u L_P=0.13u W_N=2.0u L_N=0.13u W_P_D=1.0u
+ L_P_D=0.13u W_N_D=1.0u L_N_D=0.13u n=1
*.iopin v_a
*.iopin v_b
*.iopin VDD
*.iopin VSS
*.ipin di_tg_ctrl
*.ipin di_tg_ctrl_n
XM1 v_a di_tg_ctrl v_b VSS sg13_lv_nmos w=W_N l=L_N ng=1 m=n
XM2 v_a di_tg_ctrl_n v_b VDD sg13_lv_pmos w=W_P l=L_P ng=1 m=n
XMdummy2 v_b di_tg_ctrl v_b VDD sg13_lv_pmos w=W_P_D l=L_P_D ng=1 m=n
XMdummy1 v_b di_tg_ctrl_n v_b VSS sg13_lv_nmos w=W_N_D l=L_N_D ng=1 m=n
.ends


* expanding   symbol:  inverter/inverter_lv.sym # of pins=4
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/inverter/inverter_lv.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/inverter/inverter_lv.sch
.subckt inverter_lv VDD vin vout VSS  W_P=3.0u L_P=0.13u W_N=1.0u L_N=0.13u n=1
*.ipin vin
*.iopin VDD
*.iopin VSS
*.opin vout
XM1 vout vin VDD VDD sg13_lv_pmos w=W_P l=L_P ng=1 m=n
XM2 vout vin VSS VSS sg13_lv_nmos w=W_N l=L_N ng=1 m=n
.ends


* expanding   symbol:  comparator/NOR_gate/NOR_gate.sym # of pins=5
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/comparator/NOR_gate/NOR_gate.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/comparator/NOR_gate/NOR_gate.sch
.subckt NOR_gate VDD C A B VSS  W_P=1.0u L_P=0.13u W_N=0.5u L_N=0.13u
*.iopin VDD
*.opin C
*.iopin VSS
*.ipin A
*.ipin B
XM1 C A VSS VSS sg13_lv_nmos w=W_N l=L_N ng=1 m=1
XM2 C B VSS VSS sg13_lv_nmos w=W_N l=L_N ng=1 m=1
XM3 C B net1 VDD sg13_lv_pmos w=W_P l=L_P ng=1 m=1
XM4 net1 A VDD VDD sg13_lv_pmos w=W_P l=L_P ng=1 m=1
XM5 C A net2 VDD sg13_lv_pmos w=W_P l=L_P ng=1 m=1
XM6 net2 B VDD VDD sg13_lv_pmos w=W_P l=L_P ng=1 m=1
.ends


* expanding   symbol:  transmission_gate/transmission_gate_lv_wo_dummy.sym # of pins=6
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/transmission_gate/transmission_gate_lv_wo_dummy.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/transmission_gate/transmission_gate_lv_wo_dummy.sch
.subckt transmission_gate_lv_wo_dummy VDD di_tg_ctrl VSS v_b v_a di_tg_ctrl_n  W_P=1.0u L_P=0.13u W_N=1.0u L_N=0.13u
*.iopin v_a
*.iopin v_b
*.iopin VDD
*.iopin VSS
*.ipin di_tg_ctrl
*.ipin di_tg_ctrl_n
XM1 v_a di_tg_ctrl v_b VSS sg13_lv_nmos w=W_N l=L_N ng=1 m=1
XM2 v_a di_tg_ctrl_n v_b VDD sg13_lv_pmos w=W_P l=L_P ng=1 m=1
.ends

.GLOBAL GND
**** begin user architecture code
.MODEL SW1 SW
+ VT=0.9 VH=0.01
+ RON=10 ROFF=1G
**** end user architecture code
.end
