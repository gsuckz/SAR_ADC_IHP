** sch_path: /foss/designs/SAR_ADC_IHP/xschem/comparator/NOR_gate/testbenches/NOR_gate_tb_tran.sch
**.subckt NOR_gate_tb_tran
VDD VDD GND 1.5
Vb b GND pulse(0, 1.5, 0.5n, 100p, 100p, 1n, 2n)
Va a GND pulse(0, 1.5, 0, 100p, 100p, 1n, 2n)
C1 c GND 1f m=1
R1 c GND 100Meg m=1
x1 VDD c a b GND NOR_gate W_P=1.0u L_P=0.13u W_N=0.5u L_N=0.13u
**** begin user architecture code

.lib cornerMOSlv.lib mos_tt
.lib cornerRES.lib res_typ



.param temp=27
.options savecurrents reltol=1e-3 abstol=1e-12 gmin=1e-12
.control
save all

* Operating Point Analysis
op
remzerovec
write NOR_gate_tb_tran.raw
set appendwrite

* Transient Analysis
tran 1p 4n
write NOR_gate_tb_tran.raw

plot v(A) v(B)

plot v(C)

plot i(VDD)

*quit
.endc

**** end user architecture code
**.ends

* expanding   symbol:  comparator/NOR_gate/NOR_gate.sym # of pins=5
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/comparator/NOR_gate/NOR_gate.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/comparator/NOR_gate/NOR_gate.sch
.subckt NOR_gate VDD C A B VSS  W_P=1.0u L_P=0.13u W_N=0.5u L_N=0.13u
*.iopin VDD
*.opin C
*.iopin VSS
*.ipin A
*.ipin B
XM1 C A VSS VSS sg13_lv_nmos w=W_N l=L_N ng=1 m=1
XM2 C B VSS VSS sg13_lv_nmos w=W_N l=L_N ng=1 m=1
XM3 C B net1 VDD sg13_lv_pmos w=W_P l=L_P ng=1 m=1
XM4 net1 A VDD VDD sg13_lv_pmos w=W_P l=L_P ng=1 m=1
XM5 C A net2 VDD sg13_lv_pmos w=W_P l=L_P ng=1 m=1
XM6 net2 B VDD VDD sg13_lv_pmos w=W_P l=L_P ng=1 m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.end
