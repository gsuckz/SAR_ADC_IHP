** sch_path: /foss/designs/SAR_ADC_IHP/xschem/top_level/testbenches/atbs_top_fixed_window_tb_tran.sch
**.subckt atbs_top_fixed_window_tb_tran
VDD_DAC VDD_DAC GND 1.5
VDD_COMP VDD_COMP GND 1.5
VDD_DIG VDD_DIG GND 1.5
VDD_IO VDD_IO GND 3.3
VDD_AMP VDD_AMP GND 1.5
Vcm Vcm GND 0.75
E1 Vcm vbncn net1 GND 0.5
E2 vbncp Vcm net1 GND 0.5
E3 net1 GND vsine GND 1
x1 VDD_DIG VDD_COMP clock reset_n vtrig VDD_DAC VDD_IO GND GND vecgp VDD_IO VDD_IO VDD_IO GND uart_tx idle_led overflow_led
+ underflow_led GND VDD_AMP VDD_IO vecgn vbncp vbncn vdac_uppern vdac_lowern vdac_upperp vdac_lowerp atbs_top_fixed_window
E4 Vcm vecgn net2 GND 0.5
E5 vecgp Vcm net2 GND 0.5
E6 net2 GND vecg GND 1
vsine vsine GND sin(0.75 0.65 {1/Tsig} {Tdel})
vtrig vtrig GND pulse(0 1.5 {Tdel} 10p 10p {Tsig/2} {Tsig})
vecg vecg GND dc 0 pwl(0.0 0.5958 3.910068426197458e-06 0.5985 7.820136852394917e-06 0.5982 1.1730205278592374e-05 0.6038
+ 1.5640273704789833e-05 0.61 1.9550342130987292e-05 0.6144 2.3460410557184748e-05 0.6189 2.7370478983382207e-05 0.6204 3.1280547409579666e-05 0.6162
+ 3.519061583577712e-05 0.6119 3.9100684261974585e-05 0.6106 4.301075268817204e-05 0.6123 4.6920821114369496e-05 0.6199 5.083088954056696e-05 0.6267
+ 5.4740957966764414e-05 0.6299 5.865102639296188e-05 0.6252 6.256109481915933e-05 0.6185 6.647116324535679e-05 0.6128 7.038123167155424e-05 0.6143
+ 7.429130009775171e-05 0.6176 7.820136852394917e-05 0.6242 8.211143695014662e-05 0.6294 8.602150537634408e-05 0.6272 8.993157380254154e-05 0.6273
+ 9.384164222873899e-05 0.6275 9.775171065493646e-05 0.6317 0.00010166177908113392 0.6354 0.00010557184750733137 0.6341 0.00010948191593352883 0.6258
+ 0.00011339198435972628 0.6224 0.00011730205278592375 0.6222 0.00012121212121212121 0.6297 0.00012512218963831867 0.6381 0.00012903225806451613 0.6441
+ 0.00013294232649071358 0.649 0.00013685239491691105 0.6455 0.0001407624633431085 0.6404 0.00014467253176930596 0.6344 0.00014858260019550343 0.6317
+ 0.00015249266862170087 0.6314 0.00015640273704789834 0.6377 0.00016031280547409578 0.6415 0.00016422287390029325 0.6412 0.00016813294232649072 0.643
+ 0.00017204301075268816 0.6462 0.00017595307917888563 0.6523 0.00017986314760508307 0.6546 0.00018377321603128054 0.6538 0.00018768328445747798 0.6475
+ 0.00019159335288367545 0.6412 0.00019550342130987292 0.6387 0.00019941348973607036 0.6435 0.00020332355816226783 0.6518 0.00020723362658846528 0.6618
+ 0.00021114369501466275 0.6648 0.00021505376344086021 0.6571 0.00021896383186705766 0.6539 0.00022287390029325513 0.6536 0.00022678396871945257 0.6517
+ 0.00023069403714565004 0.6562 0.0002346041055718475 0.6624 0.00023851417399804495 0.6645 0.00024242424242424242 0.6631 0.00024633431085043986 0.6616
+ 0.00025024437927663733 0.6628 0.0002541544477028348 0.6643 0.00025806451612903227 0.6666 0.0002619745845552297 0.6705 0.00026588465298142715 0.6671
+ 0.0002697947214076246 0.6628 0.0002737047898338221 0.6546 0.00027761485826001956 0.6579 0.000281524926686217 0.6719 0.00028543499511241445 0.6801
+ 0.0002893450635386119 0.6801 0.0002932551319648094 0.6725 0.00029716520039100685 0.6671 0.00030107526881720427 0.6592 0.00030498533724340174 0.6602
+ 0.0003088954056695992 0.6663 0.0003128054740957967 0.6668 0.00031671554252199415 0.6621 0.00032062561094819156 0.653 0.00032453567937438903 0.6475
+ 0.0003284457478005865 0.6456 0.00033235581622678397 0.6458 0.00033626588465298144 0.6442 0.00034017595307917885 0.6438 0.0003440860215053763 0.6375
+ 0.0003479960899315738 0.6288 0.00035190615835777126 0.6243 0.00035581622678396873 0.6349 0.00035972629521016615 0.6464 0.0003636363636363636 0.6503
+ 0.0003675464320625611 0.6447 0.00037145650048875855 0.6388 0.00037536656891495597 0.6335 0.00037927663734115344 0.6324 0.0003831867057673509 0.6363
+ 0.0003870967741935484 0.6398 0.00039100684261974585 0.6507 0.00039491691104594326 0.661 0.00039882697947214073 0.6623 0.0004027370478983382 0.6642
+ 0.00040664711632453567 0.6686 0.00041055718475073314 0.6735 0.00041446725317693055 0.6756 0.000418377321603128 0.6714 0.0004222873900293255 0.6609
+ 0.00042619745845552296 0.6532 0.00043010752688172043 0.6527 0.00043401759530791784 0.665 0.0004379276637341153 0.6815 0.0004418377321603128 0.6887
+ 0.00044574780058651025 0.6869 0.0004496578690127077 0.6736 0.00045356793743890514 0.6629 0.0004574780058651026 0.6561 0.0004613880742913001 0.6562
+ 0.00046529814271749754 0.6592 0.000469208211143695 0.6648 0.00047311827956989243 0.6671 0.0004770283479960899 0.6606 0.00048093841642228737 0.6544
+ 0.00048484848484848484 0.651 0.0004887585532746823 0.6519 0.0004926686217008797 0.6519 0.0004965786901270772 0.6545 0.0005004887585532747 0.6524
+ 0.0005043988269794721 0.6409 0.0005083088954056696 0.6268 0.000512218963831867 0.6303 0.0005161290322580645 0.6493 0.000520039100684262 0.6638
+ 0.0005239491691104594 0.6659 0.0005278592375366569 0.6581 0.0005317693059628543 0.6451 0.0005356793743890518 0.6343 0.0005395894428152492 0.6278
+ 0.0005434995112414467 0.6257 0.0005474095796676442 0.6261 0.0005513196480938416 0.6239 0.0005552297165200391 0.6154 0.0005591397849462365 0.6105
+ 0.000563049853372434 0.6115 0.0005669599217986315 0.6197 0.0005708699902248289 0.6271 0.0005747800586510264 0.6293 0.0005786901270772238 0.6242
+ 0.0005826001955034212 0.6162 0.0005865102639296188 0.6101 0.0005904203323558162 0.616 0.0005943304007820137 0.6276 0.0005982404692082111 0.6339
+ 0.0006021505376344085 0.6337 0.0006060606060606061 0.6271 0.0006099706744868035 0.6229 0.000613880742913001 0.6247 0.0006177908113391984 0.6293
+ 0.0006217008797653958 0.637 0.0006256109481915934 0.6436 0.0006295210166177908 0.643 0.0006334310850439883 0.6449 0.0006373411534701857 0.6476
+ 0.0006412512218963831 0.65 0.0006451612903225806 0.6564 0.0006490713587487781 0.6595 0.0006529814271749756 0.6571 0.000656891495601173 0.6477
+ 0.0006608015640273704 0.6374 0.0006647116324535679 0.629 0.0006686217008797654 0.6292 0.0006725317693059629 0.6357 0.0006764418377321603 0.6455
+ 0.0006803519061583577 0.6493 0.0006842619745845552 0.6455 0.0006881720430107526 0.6424 0.0006920821114369502 0.6339 0.0006959921798631476 0.625
+ 0.000699902248289345 0.6209 0.0007038123167155425 0.6215 0.0007077223851417399 0.6246 0.0007116324535679375 0.6282 0.0007155425219941349 0.6317
+ 0.0007194525904203323 0.6381 0.0007233626588465298 0.6501 0.0007272727272727272 0.6566 0.0007311827956989248 0.6539 0.0007350928641251222 0.6482
+ 0.0007390029325513196 0.6382 0.0007429130009775171 0.6283 0.0007468230694037145 0.6334 0.0007507331378299119 0.6477 0.0007546432062561095 0.6578
+ 0.0007585532746823069 0.6583 0.0007624633431085044 0.6561 0.0007663734115347018 0.6535 0.0007702834799608992 0.6449 0.0007741935483870968 0.639
+ 0.0007781036168132942 0.6398 0.0007820136852394917 0.6485 0.0007859237536656891 0.6535 0.0007898338220918865 0.6513 0.000793743890518084 0.6483
+ 0.0007976539589442815 0.6442 0.000801564027370479 0.6384 0.0008054740957966764 0.6345 0.0008093841642228738 0.6283 0.0008132942326490713 0.6215
+ 0.0008172043010752688 0.6179 0.0008211143695014663 0.6204 0.0008250244379276637 0.6304 0.0008289345063538611 0.6402 0.0008328445747800586 0.6415
+ 0.000836754643206256 0.6331 0.0008406647116324536 0.6263 0.000844574780058651 0.6245 0.0008484848484848484 0.6254 0.0008523949169110459 0.6298
+ 0.0008563049853372433 0.632 0.0008602150537634409 0.635 0.0008641251221896383 0.6377 0.0008680351906158357 0.6337 0.0008719452590420332 0.6286
+ 0.0008758553274682306 0.6293 0.0008797653958944282 0.6387 0.0008836754643206256 0.6455 0.000887585532746823 0.6419 0.0008914956011730205 0.631
+ 0.0008954056695992179 0.6165 0.0008993157380254154 0.6051 0.0009032258064516129 0.6102 0.0009071358748778103 0.6259 0.0009110459433040078 0.6371
+ 0.0009149560117302052 0.6451 0.0009188660801564027 0.6449 0.0009227761485826002 0.642 0.0009266862170087976 0.6356 0.0009305962854349951 0.629
+ 0.0009345063538611925 0.6259 0.00093841642228739 0.6271 0.0009423264907135874 0.6295 0.0009462365591397849 0.6266 0.0009501466275659824 0.6267
+ 0.0009540566959921798 0.6312 0.0009579667644183773 0.639 0.0009618768328445747 0.6441 0.0009657869012707722 0.6462 0.0009696969696969697 0.6429
+ 0.0009736070381231671 0.6387 0.0009775171065493646 0.6335 0.000981427174975562 0.6408 0.0009853372434017594 0.6532 0.0009892473118279569 0.6535
+ 0.0009931573802541545 0.6446 0.000997067448680352 0.6334 0.0010009775171065493 0.6282 0.0010048875855327467 0.6231 0.0010087976539589442 0.6265
+ 0.0010127077223851418 0.6331 0.0010166177908113392 0.6414 0.0010205278592375366 0.6474 0.001024437927663734 0.645 0.0010283479960899314 0.639
+ 0.001032258064516129 0.632 0.0010361681329423265 0.6239 0.001040078201368524 0.6222 0.0010439882697947213 0.627 0.0010478983382209187 0.6249
+ 0.0010518084066471164 0.6219 0.0010557184750733138 0.617 0.0010596285434995112 0.6225 0.0010635386119257086 0.6306 0.001067448680351906 0.6294
+ 0.0010713587487781037 0.6244 0.001075268817204301 0.6201 0.0010791788856304985 0.6194 0.001083088954056696 0.6232 0.0010869990224828933 0.6285
+ 0.001090909090909091 0.6282 0.0010948191593352884 0.6291 0.0010987292277614858 0.6302 0.0011026392961876832 0.6277 0.0011065493646138806 0.6253
+ 0.0011104594330400782 0.6244 0.0011143695014662757 0.6257 0.001118279569892473 0.6244 0.0011221896383186705 0.6272 0.001126099706744868 0.6286
+ 0.0011300097751710655 0.6217 0.001133919843597263 0.6145 0.0011378299120234604 0.6168 0.0011417399804496578 0.6251 0.0011456500488758552 0.6334
+ 0.0011495601173020528 0.6396 0.0011534701857282502 0.6362 0.0011573802541544477 0.6278 0.001161290322580645 0.616 0.0011652003910068425 0.6127
+ 0.0011691104594330401 0.6151 0.0011730205278592375 0.6206 0.001176930596285435 0.6274 0.0011808406647116324 0.6268 0.0011847507331378298 0.6251
+ 0.0011886608015640274 0.6268 0.0011925708699902248 0.6305 0.0011964809384164222 0.6318 0.0012003910068426197 0.6323 0.001204301075268817 0.6264
+ 0.0012082111436950147 0.6211 0.0012121212121212121 0.6198 0.0012160312805474095 0.6259 0.001219941348973607 0.632 0.0012238514173998044 0.633
+ 0.001227761485826002 0.636 0.0012316715542521994 0.6335 0.0012355816226783968 0.6281 0.0012394916911045942 0.6258 0.0012434017595307917 0.6319
+ 0.0012473118279569893 0.637 0.0012512218963831867 0.6389 0.0012551319648093841 0.6384 0.0012590420332355815 0.6327 0.001262952101661779 0.6333
+ 0.0012668621700879766 0.6398 0.001270772238514174 0.6508 0.0012746823069403714 0.6614 0.0012785923753665688 0.6629 0.0012825024437927662 0.6554
+ 0.0012864125122189639 0.6487 0.0012903225806451613 0.6476 0.0012942326490713587 0.6564 0.0012981427174975561 0.6702 0.0013020527859237535 0.679
+ 0.0013059628543499512 0.6801 0.0013098729227761486 0.6732 0.001313782991202346 0.6701 0.0013176930596285434 0.6706 0.0013216031280547408 0.6722
+ 0.0013255131964809385 0.6724 0.0013294232649071359 0.6741 0.0013333333333333333 0.6714 0.0013372434017595307 0.6649 0.0013411534701857281 0.6606
+ 0.0013450635386119258 0.6595 0.0013489736070381232 0.6638 0.0013528836754643206 0.6658 0.001356793743890518 0.664 0.0013607038123167154 0.6556
+ 0.001364613880742913 0.6455 0.0013685239491691105 0.6396 0.0013724340175953079 0.6482 0.0013763440860215053 0.6591 0.0013802541544477027 0.662
+ 0.0013841642228739003 0.6594 0.0013880742913000978 0.6508 0.0013919843597262952 0.6443 0.0013958944281524926 0.6412 0.00139980449657869 0.6391
+ 0.0014037145650048876 0.64 0.001407624633431085 0.6457 0.0014115347018572825 0.6474 0.0014154447702834799 0.6436 0.0014193548387096773 0.6374
+ 0.001423264907135875 0.6343 0.0014271749755620723 0.6352 0.0014310850439882698 0.6353 0.0014349951124144672 0.6288 0.0014389051808406646 0.6168
+ 0.0014428152492668622 0.5964 0.0014467253176930596 0.5828 0.001450635386119257 0.5848 0.0014545454545454545 0.5932 0.0014584555229716519 0.5988
+ 0.0014623655913978495 0.6013 0.001466275659824047 0.5993 0.0014701857282502443 0.5925 0.0014740957966764417 0.5869 0.0014780058651026392 0.5871
+ 0.0014819159335288368 0.5902 0.0014858260019550342 0.5972 0.0014897360703812316 0.6052 0.001493646138807429 0.6056 0.0014975562072336265 0.6105
+ 0.0015014662756598239 0.6175 0.0015053763440860215 0.6238 0.001509286412512219 0.6242 0.0015131964809384163 0.6232 0.0015171065493646137 0.6199
+ 0.0015210166177908112 0.6155 0.0015249266862170088 0.6119 0.0015288367546432062 0.6176 0.0015327468230694036 0.6299 0.001536656891495601 0.6393
+ 0.0015405669599217985 0.6419 0.001544477028347996 0.6374 0.0015483870967741935 0.6291 0.001552297165200391 0.6229 0.0015562072336265883 0.6219
+ 0.0015601173020527857 0.625 0.0015640273704789834 0.6286 0.0015679374389051808 0.6267 0.0015718475073313782 0.6183 0.0015757575757575756 0.6137
+ 0.001579667644183773 0.6122 0.0015835777126099707 0.6148 0.001587487781036168 0.6175 0.0015913978494623655 0.6181 0.001595307917888563 0.6126
+ 0.0015992179863147603 0.6028 0.001603128054740958 0.596 0.0016070381231671554 0.6044 0.0016109481915933528 0.6182 0.0016148582600195502 0.6263
+ 0.0016187683284457476 0.6232 0.0016226783968719453 0.6123 0.0016265884652981427 0.6041 0.00163049853372434 0.5979 0.0016344086021505375 0.5952
+ 0.001638318670576735 0.5965 0.0016422287390029325 0.6022 0.00164613880742913 0.6069 0.0016500488758553274 0.6035 0.0016539589442815248 0.603
+ 0.0016578690127077222 0.6032 0.0016617790811339198 0.6091 0.0016656891495601173 0.6148 0.0016695992179863147 0.6158 0.001673509286412512 0.6102
+ 0.0016774193548387095 0.599 0.0016813294232649071 0.5905 0.0016852394916911045 0.5946 0.001689149560117302 0.6083 0.0016930596285434994 0.6121
+ 0.0016969696969696968 0.6133 0.0017008797653958944 0.6071 0.0017047898338220918 0.5998 0.0017086999022482893 0.5943 0.0017126099706744867 0.5917
+ 0.001716520039100684 0.5903 0.0017204301075268817 0.5931 0.0017243401759530791 0.5958 0.0017282502443792765 0.5931 0.001732160312805474 0.5892
+ 0.0017360703812316714 0.5865 0.001739980449657869 0.5906 0.0017438905180840664 0.593 0.0017478005865102638 0.5958 0.0017517106549364613 0.5971
+ 0.0017556207233626587 0.592 0.0017595307917888563 0.5844 0.0017634408602150537 0.5882 0.0017673509286412511 0.5988 0.0017712609970674485 0.6044
+ 0.001775171065493646 0.6045 0.0017790811339198436 0.6 0.001782991202346041 0.5917 0.0017869012707722384 0.5876 0.0017908113391984358 0.5904
+ 0.0017947214076246333 0.5996 0.0017986314760508309 0.6059 0.0018025415444770283 0.6095 0.0018064516129032257 0.6109 0.0018103616813294231 0.6095
+ 0.0018142717497556205 0.6109 0.0018181818181818182 0.6174 0.0018220918866080156 0.6238 0.001826001955034213 0.6278 0.0018299120234604104 0.6264
+ 0.0018338220918866078 0.6177 0.0018377321603128055 0.6093 0.0018416422287390029 0.6156 0.0018455522971652003 0.6254 0.0018494623655913977 0.6305
+ 0.0018533724340175951 0.6326 0.0018572825024437928 0.6278 0.0018611925708699902 0.6259 0.0018651026392961876 0.6247 0.001869012707722385 0.6251
+ 0.0018729227761485824 0.629 0.00187683284457478 0.6279 0.0018807429130009775 0.6217 0.0018846529814271749 0.6134 0.0018885630498533723 0.6091
+ 0.0018924731182795697 0.6093 0.0018963831867057673 0.6123 0.0019002932551319648 0.6172 0.0019042033235581622 0.6183 0.0019081133919843596 0.6119
+ 0.001912023460410557 0.6026 0.0019159335288367546 0.5924 0.001919843597262952 0.5961 0.0019237536656891495 0.6095 0.0019276637341153469 0.6152
+ 0.0019315738025415443 0.6082 0.001935483870967742 0.5974 0.0019393939393939393 0.5894 0.0019433040078201368 0.5836 0.0019472140762463342 0.5864
+ 0.0019511241446725316 0.5916 0.0019550342130987292 0.5981 0.0019589442815249264 0.5983 0.001962854349951124 0.592 0.0019667644183773217 0.58
+ 0.001970674486803519 0.5702 0.0019745845552297165 0.5708 0.0019784946236559137 0.5752 0.0019824046920821113 0.5777 0.001986314760508309 0.578
+ 0.001990224828934506 0.5793 0.001994134897360704 0.5826 0.001998044965786901 0.5978 0.0020019550342130986 0.6213 0.0020058651026392963 0.6388
+ 0.0020097751710654935 0.6554 0.002013685239491691 0.6703 0.0020175953079178883 0.6918 0.002021505376344086 0.7181 0.0020254154447702836 0.7519
+ 0.0020293255131964808 0.7929 0.0020332355816226784 0.8382 0.0020371456500488756 0.8855 0.0020410557184750732 0.9325 0.002044965786901271 0.9836
+ 0.002048875855327468 1.0344 0.0020527859237536657 1.0885 0.002056695992179863 1.1466 0.0020606060606060605 1.2035 0.002064516129032258 1.2532
+ 0.0020684261974584553 1.3 0.002072336265884653 1.2942 0.00207624633431085 1.2885 0.002080156402737048 1.2826 0.0020840664711632454 1.2769
+ 0.0020879765395894426 1.2714 0.0020918866080156403 1.2668 0.0020957966764418375 1.2598 0.002099706744868035 1.2536 0.0021036168132942327 1.2482
+ 0.00210752688172043 1.2423 0.0021114369501466276 1.2365 0.0021153470185728248 1.231 0.0021192570869990224 1.2252 0.00212316715542522 1.2196
+ 0.0021270772238514172 1.2133 0.002130987292277615 1.1967 0.002134897360703812 1.1296 0.0021388074291300097 1.0419 0.0021427174975562073 0.9281
+ 0.0021466275659824045 0.8036 0.002150537634408602 0.6811 0.0021544477028347993 0.5654 0.002158357771260997 0.4556 0.0021622678396871946 0.3608
+ 0.002166177908113392 0.2826 0.0021700879765395894 0.217 0.0021739980449657866 0.1684 0.0021779081133919843 0.1376 0.002181818181818182 0.1154
+ 0.002185728250244379 0.1 0.0021896383186705767 0.1009 0.002193548387096774 0.1122 0.0021974584555229716 0.1309 0.002201368523949169 0.159
+ 0.0022052785923753664 0.1921 0.002209188660801564 0.2272 0.0022130987292277612 0.2652 0.002217008797653959 0.2953 0.0022209188660801565 0.3131
+ 0.0022248289345063537 0.3249 0.0022287390029325513 0.3361 0.0022326490713587485 0.3577 0.002236559139784946 0.382 0.0022404692082111438 0.3989
+ 0.002244379276637341 0.4072 0.0022482893450635386 0.4052 0.002252199413489736 0.4011 0.0022561094819159334 0.3957 0.002260019550342131 0.3998
+ 0.0022639296187683283 0.4047 0.002267839687194526 0.4115 0.002271749755620723 0.4171 0.0022756598240469207 0.4189 0.0022795698924731184 0.4211
+ 0.0022834799608993156 0.4295 0.002287390029325513 0.4436 0.0022913000977517104 0.453 0.002295210166177908 0.4584 0.0022991202346041057 0.4591
+ 0.002303030303030303 0.4579 0.0023069403714565005 0.4602 0.0023108504398826977 0.4714 0.0023147605083088953 0.4834 0.002318670576735093 0.487
+ 0.00232258064516129 0.4845 0.0023264907135874878 0.4786 0.002330400782013685 0.4672 0.0023343108504398826 0.4578 0.0023382209188660802 0.4515
+ 0.0023421309872922774 0.4524 0.002346041055718475 0.4611 0.0023499511241446723 0.4644 0.00235386119257087 0.4609 0.0023577712609970675 0.4619
+ 0.0023616813294232647 0.4655 0.0023655913978494624 0.4743 0.0023695014662756596 0.4811 0.002373411534701857 0.4826 0.002377321603128055 0.4771
+ 0.002381231671554252 0.4694 0.0023851417399804497 0.4687 0.002389051808406647 0.478 0.0023929618768328445 0.4897 0.002396871945259042 0.4957
+ 0.0024007820136852393 0.5 0.002404692082111437 0.4979 0.002408602150537634 0.4968 0.0024125122189638318 0.4965 0.0024164222873900294 0.5002
+ 0.0024203323558162266 0.5095 0.0024242424242424242 0.5165 0.0024281524926686214 0.5223 0.002432062561094819 0.5205 0.0024359726295210167 0.5186
+ 0.002439882697947214 0.5205 0.0024437927663734115 0.5281 0.0024477028347996087 0.5415 0.0024516129032258064 0.5447 0.002455522971652004 0.5397
+ 0.002459433040078201 0.5315 0.002463343108504399 0.5274 0.002467253176930596 0.535 0.0024711632453567937 0.5484 0.0024750733137829913 0.5567
+ 0.0024789833822091885 0.5636 0.002482893450635386 0.5627 0.0024868035190615833 0.5603 0.002490713587487781 0.5545 0.0024946236559139786 0.5528
+ 0.0024985337243401758 0.5518 0.0025024437927663734 0.553 0.0025063538611925706 0.5516 0.0025102639296187682 0.5499 0.002514173998044966 0.5449
+ 0.002518084066471163 0.5471 0.0025219941348973607 0.5603 0.002525904203323558 0.5685 0.0025298142717497555 0.572 0.002533724340175953 0.5676
+ 0.0025376344086021504 0.5602 0.002541544477028348 0.5534 0.002545454545454545 0.5604 0.002549364613880743 0.5731 0.0025532746823069405 0.5841
+ 0.0025571847507331377 0.5875 0.0025610948191593353 0.5869 0.0025650048875855325 0.5827 0.00256891495601173 0.5792 0.0025728250244379277 0.5812
+ 0.002576735092864125 0.5859 0.0025806451612903226 0.5908 0.0025845552297165198 0.5914 0.0025884652981427174 0.5866 0.002592375366568915 0.5871
+ 0.0025962854349951122 0.593 0.00260019550342131 0.5996 0.002604105571847507 0.6003 0.0026080156402737047 0.5944 0.0026119257086999023 0.5892
+ 0.0026158357771260995 0.5891 0.002619745845552297 0.5901 0.0026236559139784944 0.5936 0.002627565982404692 0.6017 0.0026314760508308896 0.6066
+ 0.002635386119257087 0.6024 0.0026392961876832845 0.5985 0.0026432062561094817 0.5996 0.0026471163245356793 0.5982 0.002651026392961877 0.5962
+ 0.002654936461388074 0.5969 0.0026588465298142717 0.6024 0.002662756598240469 0.6041 0.0026666666666666666 0.6056 0.002670576735092864 0.6091
+ 0.0026744868035190614 0.6126 0.002678396871945259 0.6169 0.0026823069403714562 0.6229 0.002686217008797654 0.6264 0.0026901270772238515 0.6181
+ 0.0026940371456500487 0.6077 0.0026979472140762463 0.6017 0.0027018572825024435 0.6124 0.002705767350928641 0.6275 0.002709677419354839 0.6336
+ 0.002713587487781036 0.6293 0.0027174975562072336 0.619 0.002721407624633431 0.6046 0.0027253176930596285 0.5948 0.002729227761485826 0.5948
+ 0.0027331378299120233 0.5995 0.002737047898338221 0.5994 0.002740957966764418 0.595 0.0027448680351906157 0.5861 0.0027487781036168134 0.5802
+ 0.0027526881720430106 0.5825 0.002756598240469208 0.5913 0.0027605083088954054 0.6001 0.002764418377321603 0.6049 0.0027683284457478007 0.6012
+ 0.002772238514173998 0.5907 0.0027761485826001955 0.585 0.0027800586510263927 0.5939 0.0027839687194525903 0.607 0.002787878787878788 0.6169
+ 0.002791788856304985 0.625 0.002795698924731183 0.6239 0.00279960899315738 0.6239 0.0028035190615835776 0.621 0.0028074291300097753 0.624
+ 0.0028113391984359725 0.6299 0.00281524926686217 0.6359 0.0028191593352883673 0.6377 0.002823069403714565 0.6335 0.0028269794721407625 0.6341
+ 0.0028308895405669597 0.6396 0.0028347996089931574 0.6458 0.0028387096774193546 0.6499 0.002842619745845552 0.6522 0.00284652981427175 0.6458
+ 0.002850439882697947 0.6395 0.0028543499511241447 0.6349 0.002858260019550342 0.6389 0.0028621700879765395 0.6482 0.002866080156402737 0.6495
+ 0.0028699902248289343 0.6445 0.002873900293255132 0.6378 0.002877810361681329 0.6328 0.002881720430107527 0.6295 0.0028856304985337244 0.6306
+ 0.0028895405669599216 0.6367 0.0028934506353861193 0.6514 0.0028973607038123165 0.6632 0.002901270772238514 0.6617 0.0029051808406647117 0.6624
+ 0.002909090909090909 0.6643 0.0029130009775171065 0.6646 0.0029169110459433037 0.6642 0.0029208211143695014 0.6612 0.002924731182795699 0.6518
+ 0.002928641251221896 0.6433 0.002932551319648094 0.6426 0.002936461388074291 0.6522 0.0029403714565004887 0.6656 0.0029442815249266863 0.6728
+ 0.0029481915933528835 0.6738 0.002952101661779081 0.6692 0.0029560117302052783 0.666 0.002959921798631476 0.667 0.0029638318670576736 0.6666
+ 0.002967741935483871 0.6644 0.0029716520039100684 0.6657 0.0029755620723362656 0.6638 0.0029794721407624633 0.6568 0.002983382209188661 0.6551
+ 0.002987292277614858 0.6566 0.0029912023460410557 0.6631 0.002995112414467253 0.6689 0.0029990224828934505 0.6677 0.0030029325513196477 0.662
+ 0.0030068426197458454 0.6549 0.003010752688172043 0.6551 0.00301466275659824 0.6691 0.003018572825024438 0.6819 0.003022482893450635 0.6912
+ 0.0030263929618768327 0.695 0.0030303030303030303 0.6932 0.0030342130987292275 0.6952 0.003038123167155425 0.7034 0.0030420332355816223 0.7138
+ 0.00304594330400782 0.7209 0.0030498533724340176 0.7327 0.003053763440860215 0.7376 0.0030576735092864124 0.7351 0.0030615835777126096 0.7336
+ 0.0030654936461388073 0.7328 0.003069403714565005 0.7369 0.003073313782991202 0.7404 0.0030772238514173997 0.7446 0.003081133919843597 0.7451
+ 0.0030850439882697945 0.7433 0.003088954056695992 0.743 0.0030928641251221894 0.7505 0.003096774193548387 0.7563 0.003100684261974584 0.7588
+ 0.003104594330400782 0.7581 0.0031085043988269795 0.7551 0.0031124144672531767 0.7517 0.0031163245356793743 0.7522 0.0031202346041055715 0.7564
+ 0.003124144672531769 0.7643 0.0031280547409579668 0.7735 0.003131964809384164 0.7788 0.0031358748778103616 0.7806 0.003139784946236559 0.7857
+ 0.0031436950146627564 0.7898 0.003147605083088954 0.7975 0.0031515151515151513 0.8073 0.003155425219941349 0.8131 0.003159335288367546 0.816
+ 0.0031632453567937437 0.8181 0.0031671554252199413 0.8195 0.0031710654936461385 0.8293 0.003174975562072336 0.8431 0.0031788856304985334 0.8512
+ 0.003182795698924731 0.8559 0.0031867057673509286 0.8577 0.003190615835777126 0.8607 0.0031945259042033235 0.8584 0.0031984359726295207 0.8553
+ 0.0032023460410557183 0.8529 0.003206256109481916 0.849 0.003210166177908113 0.8428 0.0032140762463343108 0.8393 0.003217986314760508 0.8444
+ 0.0032218963831867056 0.8496 0.0032258064516129032 0.8541 0.0032297165200391004 0.8575 0.003233626588465298 0.8566 0.0032375366568914953 0.8492
+ 0.003241446725317693 0.8411 0.0032453567937438905 0.8339 0.0032492668621700877 0.8355 0.0032531769305962853 0.8438 0.0032570869990224825 0.849
+ 0.00326099706744868 0.8448 0.003264907135874878 0.8321 0.003268817204301075 0.8248 0.0032727272727272726 0.8203 0.00327663734115347 0.8166
+ 0.0032805474095796675 0.8224 0.003284457478005865 0.8301 0.0032883675464320623 0.8385 0.00329227761485826 0.8371 0.003296187683284457 0.8262
+ 0.0033000977517106548 0.8151 0.0033040078201368524 0.8133 0.0033079178885630496 0.8143 0.0033118279569892472 0.8109 0.0033157380254154444 0.8008
+ 0.003319648093841642 0.7874 0.0033235581622678397 0.7754 0.003327468230694037 0.7759 0.0033313782991202345 0.7809 0.0033352883675464317 0.7835
+ 0.0033391984359726293 0.7746 0.003343108504398827 0.7588 0.003347018572825024 0.75 0.003350928641251222 0.7429 0.003354838709677419 0.7373
+ 0.0033587487781036166 0.7301 0.0033626588465298143 0.727 0.0033665689149560115 0.7161 0.003370478983382209 0.696 0.0033743890518084063 0.6794
+ 0.003378299120234604 0.6727 0.0033822091886608016 0.6671 0.0033861192570869988 0.6623 0.0033900293255131964 0.6511 0.0033939393939393936 0.6306
+ 0.0033978494623655912 0.6095 0.003401759530791789 0.5925 0.003405669599217986 0.5872 0.0034095796676441837 0.5844 0.003413489736070381 0.5781
+ 0.0034173998044965785 0.5696 0.003421309872922776 0.5558 0.0034252199413489733 0.541 0.003429130009775171 0.5191 0.003433040078201368 0.5036
+ 0.003436950146627566 0.4921 0.0034408602150537634 0.4852 0.0034447702834799606 0.4715 0.0034486803519061583 0.4564 0.0034525904203323555 0.4464
+ 0.003456500488758553 0.4411 0.0034604105571847507 0.4438 0.003464320625610948 0.4418 0.0034682306940371456 0.4314 0.0034721407624633428 0.4168
+ 0.0034760508308895404 0.4047 0.003479960899315738 0.3946 0.0034838709677419352 0.3934 0.003487781036168133 0.3956 0.00349169110459433 0.3906
+ 0.0034956011730205277 0.3816 0.0034995112414467253 0.3725 0.0035034213098729225 0.3634 0.00350733137829912 0.3497 0.0035112414467253173 0.3389
+ 0.003515151515151515 0.3377 0.0035190615835777126 0.3388 0.00352297165200391 0.3349 0.0035268817204301074 0.328 0.0035307917888563046 0.3205
+ 0.0035347018572825023 0.3179 0.0035386119257087 0.3206 0.003542521994134897 0.3233 0.0035464320625610947 0.3216 0.003550342130987292 0.3157
+ 0.0035542521994134896 0.3059 0.003558162267839687 0.2951 0.0035620723362658844 0.2939 0.003565982404692082 0.3011 0.0035698924731182792 0.3006
+ 0.003573802541544477 0.2988 0.0035777126099706745 0.2972 0.0035816226783968717 0.295 0.0035855327468230693 0.2941 0.0035894428152492665 0.2993
+ 0.003593352883675464 0.3056 0.0035972629521016618 0.3162 0.003601173020527859 0.3249 0.0036050830889540566 0.3257 0.003608993157380254 0.3269
+ 0.0036129032258064514 0.3268 0.003616813294232649 0.3276 0.0036207233626588463 0.331 0.003624633431085044 0.3277 0.003628543499511241 0.3258
+ 0.0036324535679374387 0.3218 0.0036363636363636364 0.3131 0.0036402737047898336 0.3214 0.003644183773216031 0.3389 0.0036480938416422284 0.3469
+ 0.003652003910068426 0.3501 0.0036559139784946237 0.3423 0.003659824046920821 0.3349 0.0036637341153470185 0.3292 0.0036676441837732157 0.3288
+ 0.0036715542521994133 0.3339 0.003675464320625611 0.3474 0.003679374389051808 0.3572 0.0036832844574780058 0.3568 0.003687194525904203 0.3557
+ 0.0036911045943304006 0.3541 0.0036950146627565982 0.3578 0.0036989247311827954 0.3649 0.003702834799608993 0.3709 0.0037067448680351903 0.3746
+ 0.003710654936461388 0.3741 0.0037145650048875855 0.3726 0.0037184750733137827 0.3857 0.0037223851417399804 0.4015 0.0037262952101661776 0.4087
+ 0.003730205278592375 0.4071 0.003734115347018573 0.4036 0.00373802541544477 0.4005 0.0037419354838709677 0.4027 0.003745845552297165 0.4112
+ 0.0037497556207233625 0.4201 0.00375366568914956 0.4278 0.0037575757575757573 0.4325 0.003761485826001955 0.433 0.003765395894428152 0.4363
+ 0.0037693059628543498 0.4351 0.0037732160312805474 0.4349 0.0037771260997067446 0.4367 0.0037810361681329422 0.4386 0.0037849462365591394 0.4376
+ 0.003788856304985337 0.4372 0.0037927663734115347 0.4351 0.003796676441837732 0.4419 0.0038005865102639295 0.4512 0.0038044965786901267 0.4559
+ 0.0038084066471163244 0.457 0.003812316715542522 0.4584 0.003816226783968719 0.4638 0.003820136852394917 0.469 0.003824046920821114 0.4758
+ 0.0038279569892473117 0.4785 0.0038318670576735093 0.4824 0.0038357771260997065 0.4866 0.003839687194525904 0.4862 0.0038435972629521013 0.4888
+ 0.003847507331378299 0.4946 0.0038514173998044966 0.5018 0.0038553274682306938 0.511 0.0038592375366568914 0.5156 0.0038631476050830886 0.516
+ 0.0038670576735092862 0.5103 0.003870967741935484 0.5061 0.003874877810361681 0.5146 0.0038787878787878787 0.5265 0.003882697947214076 0.5318
+ 0.0038866080156402735 0.5323 0.003890518084066471 0.5304 0.0038944281524926684 0.5326 0.003898338220918866 0.5327 0.003902248289345063 0.5336
+ 0.003906158357771261 0.5339 0.0039100684261974585 0.5347 0.003913978494623656 0.5356 0.003917888563049853 0.5347 0.003921798631476051 0.5355
+ 0.003925708699902248 0.5417 0.003929618768328445 0.5518 0.003933528836754643 0.5575 0.003937438905180841 0.5562 0.003941348973607038 0.5498
+ 0.003945259042033236 0.5394 0.003949169110459433 0.5324 0.00395307917888563 0.5382 0.003956989247311827 0.5497 0.0039608993157380255 0.5578
+ 0.003964809384164223 0.5558 0.00396871945259042 0.554 0.003972629521016618 0.5549 0.003976539589442815 0.5578 0.003980449657869012 0.5618
+ 0.00398435972629521 0.5665 0.003988269794721408 0.5743 0.003992179863147605 0.5782 0.003996089931573802 0.5752 0.004 0.5699 )
vrst reset_n GND pulse(1.5 0 {2/fclk} 10p 10p {2/fclk} 1 1)
vclk clock GND pulse(0 1.5 0 10p 10p {0.5/fclk} {1/fclk})
**** begin user architecture code



* Gate-Level Analog Mixed Signal Simulation (.xspice)
.include /foss/designs/SG13G2_ATBS-ADC-main/xspice/atbs_core_fixed_window_board/atbs_core_fixed_window_board.xspice
.param temp=27
.param fclk=8000000
.csparam fclk=fclk
*.param Tsig=20m
*.param Tdel=20m
.param Tsig=200u
.param Tdel=100u
.csparam Tsig=Tsig
.csparam Tdel=Tdel
.options savecurrents method=gear reltol=1e-2 abstol=1e-12 gmin=1e-12 rshunt=1e12
.control

* save all
save vecg vecgp vecgn vbnc vbncp vbncn vtrig clock reset_n uart_tx idle_led overflow_led underflow_led vdac_upperp vdac_uppern vdac_lowerp vdac_lowern
save x1.Vcm x1.voutp_amp x1.voutn_amp x1.voutp_switch x1.voutn_switch
save x1.spike x1.bio_amp_en x1.en_cap_1 x1.en_cap_2 x1.en_cap_3 x1.spdt_ctrl
save x1.phi_vcm_generator_1 x1.phi_vcm_generator_2 x1.phi_bias_1 x1.phi_bias_2 x1.phi_cmfb_1 x1.phi_cmfb_2 x1.phi_R_1 x1.phi_R_2
save x1.phi_comp x1.vcomp_upper x1.vcomp_lower x1.phi_dac_upper x1.dac_D0_upper x1.dac_D1_upper x1.dac_D2_upper x1.dac_D3_upper x1.phi_dac_lower x1.dac_D0_lower x1.dac_D1_lower x1.dac_D2_lower x1.dac_D3_lower

* Transient Analysis
let tstep = 1/fclk
let tstop = Tdel + 4*Tsig
tran $&tstep $&tstop
write atbs_top_fixed_window_tb_tran.raw

* Plotting Data
let vdac_upper = vdac_upperp - vdac_uppern
let vdac_lower = vdac_lowerp - vdac_lowern
plot v(vecg) v(vsine) v(vtrig) v(vdac_upper) v(vdac_lower)

* Calculate Energy / Conversion (ToDo for all VDDs and add together in the end)
* i_int in As
* energy_conv in Ws = J
* let N = 1
* let t_conv = 1/fclk
* meas tran i_int INTEG i(VDD) from=0p to=t_conv
* let energy_conv = 1.5 * i_int / N

* let energy_conv_pico = energy_conv * 1e12
* echo Energy / Conversion $&energy_conv_pico pJ/conv

* Calculate Power Consumption (ToDo)
* let power = energy_conv / t_conv * 1e6
* echo Power Consumption $&power uW

* Writing Data
set wr_singlescale
set wr_vecnames
wrdata /foss/designs/SG13G2_ATBS-ADC-main/python/plot_simulations/data/atbs_top_fixed_window_tb_tran.txt v(vecg) v(vsine) v(vdac_upper) v(vdac_lower)
wrdata /foss/designs/SG13G2_ATBS-ADC-main/python/reconstruction/data/atbs_top_fixed_window_tb_tran_uart.txt v(clock) v(uart_tx)
set appendwrite

.endc




.lib cornerMOSlv.lib mos_tt
.lib cornerMOShv.lib mos_tt
.lib cornerRES.lib res_typ
.include sg13g2_esd.lib


**** end user architecture code
**.ends

* expanding   symbol:  top_level/atbs_top_fixed_window.sym # of pins=28
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/top_level/atbs_top_fixed_window.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/top_level/atbs_top_fixed_window.sch
.subckt atbs_top_fixed_window VDD_DIG VDD_COMP di_clock di_reset_n di_trigger_start_sampling VDD_DAC di_trigger_start_mode
+ di_adaptive_mode di_control_mode vecgp di_signal_select_in di_enable di_select_tbs_delta_steps di_uart_rx do_uart_tx do_idle_led do_overflow_led
+ do_underflow_led VSS VDD_AMP VDD_IO vecgn vbncp vbncn vdac_uppern vdac_lowern vdac_upperp vdac_lowerp
*.iopin VDD_DIG
*.iopin VSS
*.iopin VDD_COMP
*.ipin vecgp
*.ipin di_clock
*.ipin di_reset_n
*.iopin VDD_DAC
*.ipin di_uart_rx
*.opin do_uart_tx
*.ipin di_trigger_start_sampling
*.ipin di_trigger_start_mode
*.ipin di_adaptive_mode
*.ipin di_control_mode
*.ipin di_signal_select_in
*.ipin di_enable
*.ipin di_select_tbs_delta_steps
*.opin do_idle_led
*.opin do_overflow_led
*.opin do_underflow_led
*.opin vdac_upperp
*.opin vdac_lowern
*.iopin VDD_AMP
*.ipin vecgn
*.ipin vbncp
*.ipin vbncn
*.iopin VDD_IO
*.opin vdac_uppern
*.opin vdac_lowerp
x1 phi_bias_2_buf phi_bias_1_buf phi_R_2_buf phi_R_1_buf en_cap_3_buf en_cap_1_buf en_cap_2_buf phi_cmfb_2_buf phi_cmfb_1_buf
+ voutp_amp bio_amp_en_buf net1 Vcm voutn_amp net2 VDD_AMP VSS bio_amplifier
x2 VDD_DIG spdt_ctrl_buf VSS voutn_switch net4 voutn_amp spdt_switch W_P_TG=3.0u L_P_TG=0.13u W_N_TG=1.0u L_N_TG=0.13u
x3 VDD_DIG spdt_ctrl_buf VSS voutp_switch net3 voutp_amp spdt_switch W_P_TG=3.0u L_P_TG=0.13u W_N_TG=1.0u L_N_TG=0.13u
x4 VDD_COMP vdac_upperp vcomp_upper vdac_uppern phi_comp_buf VSS DT_comparator
x5 VDD_COMP vdac_lowerp vcomp_lower vdac_lowern phi_comp_buf VSS DT_comparator
x30 VDD_DIG VSS adaptive_mode bio_amp_en clock vcomp_lower vcomp_upper control_mode dac_D0_lower dac_D1_lower dac_D2_lower
+ dac_D3_lower dac_D0_upper dac_D1_upper dac_D2_upper dac_D3_upper enable idle_led overflow_led phi_bias_1 phi_bias_2 phi_cmfb_1 phi_cmfb_2
+ phi_comp phi_dac_lower phi_dac_upper phi_R_1 phi_R_2 phi_vcm_generator_1 phi_vcm_generator_2 reset_n en_cap_1 en_cap_2 en_cap_3 spdt_ctrl
+ select_tbs_delta_steps signal_select_in spike trigger_start_mode trigger_start_sampling uart_rx uart_tx underflow_led atbs_core_fixed_window_board
x32 VDD_DIG phi_vcm_generator_2_buf phi_vcm_generator_1_buf Vcm VSS vcm_generator C_VCM=1p W_P_VCM=1.0u L_P_VCM=0.13u W_N_VCM=1.0u
+ L_N_VCM=0.13u
x31 VDD_DAC voutp_switch vdac_upperp vdac_uppern voutn_switch dac_D0_lower_buf dac_D1_lower_buf dac_D2_lower_buf dac_D3_lower_buf
+ VSS VDD_DAC Vcm vdac_lowerp vdac_lowern phi_dac_lower_buf dac_D0_upper_buf dac_D1_upper_buf dac_D2_upper_buf dac_D3_upper_buf
+ phi_dac_upper_buf dac W_P_SPDT=1.0u L_P_SPDT=0.13u W_N_SPDT=1.0u L_N_SPDT=0.13u C2=1024f Cu=8f Cucomp=8.1f
x6 VDD_IO di_clock di_control_mode clock control_mode VSS di_reset_n reset_n di_signal_select_in signal_select_in enable
+ trigger_start_sampling di_trigger_start_sampling di_enable select_tbs_delta_steps di_select_tbs_delta_steps trigger_start_mode di_trigger_start_mode
+ di_adaptive_mode uart_rx adaptive_mode di_uart_rx VDD_DIG input_hardware
x7 uart_tx do_uart_tx do_idle_led idle_led do_overflow_led overflow_led underflow_led do_underflow_led VDD_IO VSS VDD_DIG
+ output_hardware
x8 VDD_AMP vecgp net1 VSS esd_protection
x9 VDD_AMP vecgn net2 VSS esd_protection
x10 VDD_DIG phi_dac_lower phi_bias_1_buf phi_dac_upper phi_cmfb_1 phi_dac_lower_buf phi_cmfb_1_buf phi_bias_1 phi_dac_upper_buf
+ VSS dac_D0_lower dac_D0_lower_buf phi_cmfb_2 phi_bias_2_buf phi_bias_2 dac_D0_upper dac_D0_upper_buf phi_cmfb_2_buf dac_D1_upper
+ phi_R_1_buf phi_R_1 en_cap_1_buf dac_D1_lower_buf dac_D1_upper_buf dac_D1_lower en_cap_1 dac_D2_upper phi_R_2_buf phi_R_2 en_cap_2_buf
+ dac_D2_lower_buf en_cap_2 dac_D2_lower dac_D2_upper_buf bio_amp_en_buf en_cap_3_buf en_cap_3 bio_amp_en dac_D3_upper_buf dac_D3_lower_buf
+ dac_D3_lower dac_D3_upper phi_comp phi_vcm_generator_1_buf phi_vcm_generator_1 spdt_ctrl_buf spdt_ctrl phi_comp_buf phi_vcm_generator_2_buf
+ phi_vcm_generator_2 buffers
x11 VDD_AMP vbncp net3 VSS esd_protection
x12 VDD_AMP vbncn net4 VSS esd_protection
.ends


* expanding   symbol:  bio_amplifier/bio_amplifier.sym # of pins=17
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/bio_amplifier/bio_amplifier.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/bio_amplifier/bio_amplifier.sch
.subckt bio_amplifier di_phi_bias_2 di_phi_bias_1 di_phi_R_2 di_phi_R_1 di_en_cap_3 di_en_cap_1 di_en_cap_2 di_phi_cmfb_2
+ di_phi_cmfb_1 voutp di_bio_amp_en vinp Vcm voutn vinn VDD VSS
*.iopin VDD
*.iopin VSS
*.ipin di_bio_amp_en
*.ipin vinp
*.ipin vinn
*.ipin Vcm
*.opin voutp
*.opin voutn
*.ipin di_phi_cmfb_1
*.ipin di_phi_cmfb_2
*.ipin di_phi_R_1
*.ipin di_phi_R_2
*.ipin di_phi_bias_1
*.ipin di_phi_bias_2
*.ipin di_en_cap_1
*.ipin di_en_cap_2
*.ipin di_en_cap_3
x2 net1 voutn di_phi_R_2 di_phi_R_1 VDD VSS sc_fb_resistor W_P_FB=1.0u L_P_FB=0.13u W_N_FB=1.0u L_N_FB=0.13u Cs=4f
x3 net2 voutp di_phi_R_2 di_phi_R_1 VDD VSS sc_fb_resistor W_P_FB=1.0u L_P_FB=0.13u W_N_FB=1.0u L_N_FB=0.13u Cs=4f
C2a voutn net1 3.3p m=1
C2b voutp net2 3.3p m=1
x4 VDD di_en_cap_1 VSS di_en_cap_2 vinp net1 di_en_cap_3 programmable_cap_x3 W_P_PC=1.0u L_P_PC=0.13u W_N_PC=1.0u L_N_PC=0.13u
+ C1=33p C2=132p C3=165p
x5 VDD di_en_cap_1 VSS di_en_cap_2 vinn net2 di_en_cap_3 programmable_cap_x3 W_P_PC=1.0u L_P_PC=0.13u W_N_PC=1.0u L_N_PC=0.13u
+ C1=33p C2=132p C3=165p
x1 di_phi_cmfb_1 di_phi_bias_2 di_phi_bias_1 di_phi_cmfb_2 voutp voutn di_bio_amp_en net2 net1 VDD VSS Vcm amplifier_core
.ends


* expanding   symbol:  spdt_switch/spdt_switch.sym # of pins=6
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/spdt_switch/spdt_switch.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/spdt_switch/spdt_switch.sch
.subckt spdt_switch VDD di_spdt_ctrl VSS v_c v_b v_a  W_P_TG=3.0u L_P_TG=0.13u W_N_TG=1.0u L_N_TG=0.13u
*.iopin v_a
*.iopin v_b
*.iopin v_c
*.iopin VDD
*.iopin VSS
*.ipin di_spdt_ctrl
x1 VDD di_spdt_ctrl VSS v_c v_a di_spdt_ctrl_n transmission_gate_lv_wo_dummy W_P=W_P_TG L_P=L_P_TG W_N=W_N_TG L_N=L_N_TG
x2 VDD di_spdt_ctrl_n VSS v_b v_c di_spdt_ctrl transmission_gate_lv_wo_dummy W_P=W_P_TG L_P=L_P_TG W_N=W_N_TG L_N=L_N_TG
x8 VDD di_spdt_ctrl di_spdt_ctrl_n VSS inverter_lv W_P=W_P_TG L_P=L_P_TG W_N=W_N_TG L_N=L_N_TG
.ends


* expanding   symbol:  comparator/discrete_time/DT_comparator.sym # of pins=6
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/comparator/discrete_time/DT_comparator.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/comparator/discrete_time/DT_comparator.sch
.subckt DT_comparator VDD vinp vout vinn di_clk VSS
*.iopin VDD
*.opin vout
*.iopin VSS
*.ipin vinp
*.ipin vinn
*.ipin di_clk
x2 VDD voutp_comp voutp_buf VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x3 VDD voutn_comp voutn_buf VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x5 VDD di_clk net1 VSS inverter_lv W_P=1.0u L_P=0.13u W_N=1.0u L_N=0.13u
* noconn #net2
x4 VDD voutp_buf net2 VSS vout voutn_buf SR_latch W_P_SR=1.0u L_P_SR=0.13u W_N_SR=1.0u L_N_SR=0.13u
x1 net1 di_clk VDD voutp_comp vinp VSS voutn_comp vinn dynamic_biasing_comparator
.ends


* expanding   symbol:  vcm_generator/vcm_generator.sym # of pins=5
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/vcm_generator/vcm_generator.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/vcm_generator/vcm_generator.sch
.subckt vcm_generator VDD di_phi_2 di_phi_1 Vcm VSS  C_VCM=1p W_P_VCM=1.0u L_P_VCM=0.13u W_N_VCM=1.0u L_N_VCM=0.13u
*.iopin VDD
*.opin Vcm
*.iopin VSS
*.ipin di_phi_1
*.ipin di_phi_2
x1 VDD di_phi_2 VSS net1 VDD di_phi_2_n transmission_gate_lv_wo_dummy W_P=W_P_VCM L_P=L_P_VCM W_N=W_N_VCM L_N=L_N_VCM
x2 VDD di_phi_1 VSS Vcm net1 di_phi_1_n transmission_gate_lv_wo_dummy W_P=W_P_VCM L_P=L_P_VCM W_N=W_N_VCM L_N=L_N_VCM
x3 VDD di_phi_2 VSS net3 net2 di_phi_2_n transmission_gate_lv_wo_dummy W_P=W_P_VCM L_P=L_P_VCM W_N=W_N_VCM L_N=L_N_VCM
x4 VDD di_phi_1 VSS Vcm net3 di_phi_1_n transmission_gate_lv_wo_dummy W_P=W_P_VCM L_P=L_P_VCM W_N=W_N_VCM L_N=L_N_VCM
x5 VDD di_phi_1 VSS VSS net2 di_phi_1_n transmission_gate_lv_wo_dummy W_P=W_P_VCM L_P=L_P_VCM W_N=W_N_VCM L_N=L_N_VCM
x9 VDD di_phi_1 di_phi_1_n VSS inverter_lv W_P=W_P_VCM L_P=L_P_VCM W_N=W_N_VCM L_N=L_N_VCM
x8 VDD di_phi_2 di_phi_2_n VSS inverter_lv W_P=W_P_VCM L_P=L_P_VCM W_N=W_N_VCM L_N=L_N_VCM
C1 net1 net2 C_VCM m=1
C2 net3 VSS C_VCM m=1
.ends


* expanding   symbol:  dac/dac.sym # of pins=20
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/dac/dac.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/dac/dac.sch
.subckt dac VDD vinp voutp1 voutn1 vinn di_D0_2 di_D1_2 di_D2_2 di_D3_2 VSS Vref Vcm voutp2 voutn2 di_clk_2 di_D0_1 di_D1_1
+ di_D2_1 di_D3_1 di_clk_1  W_P_SPDT=1.0u L_P_SPDT=0.13u W_N_SPDT=1.0u L_N_SPDT=0.13u C2=1024f Cu=8f Cucomp=8.1f
*.opin voutp1
*.ipin di_D0_1
*.iopin VSS
*.iopin Vref
*.opin voutn1
*.ipin vinp
*.ipin vinn
*.ipin di_D1_1
*.ipin di_D2_1
*.ipin di_D3_1
*.opin voutp2
*.opin voutn2
*.iopin VDD
*.ipin Vcm
*.ipin di_clk_1
*.ipin di_D3_2
*.ipin di_D2_2
*.ipin di_D1_2
*.ipin di_D0_2
*.ipin di_clk_2
C2a vinp voutp1 C2 m=1
C2b vinn voutn1 C2 m=1
C1a net3 voutp1 Cucomp m=1
C1b net1 voutn1 Cucomp m=1
x2 VDD di_clk_1 VSS voutp1 Vcm clk_1_n transmission_gate_lv_wo_dummy W_P=1.0u L_P=0.13u W_N=1.0u L_N=0.13u
x3 VDD di_clk_1 VSS voutn1 Vcm clk_1_n transmission_gate_lv_wo_dummy W_P=1.0u L_P=0.13u W_N=1.0u L_N=0.13u
x1 VDD di_clk_1 clk_1_n VSS inverter_lv W_P=W_P_SPDT L_P=L_P_SPDT W_N=W_N_SPDT L_N=L_N_SPDT
x5 Vref VSS VSS di_D1_1 di_clk_1 VDD voutp1 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=2*Cu
x6 Vref VSS VSS di_D2_1 di_clk_1 VDD voutp1 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=4*Cu
x4 Vref VSS VSS di_D0_1 di_clk_1 VDD voutp1 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=Cu
x7 Vref VSS VSS di_D3_1 di_clk_1 VDD voutp1 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=8*Cu
x9 VSS Vref VSS di_D0_1 di_clk_1 VDD voutn1 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=Cu
x10 VSS Vref VSS di_D1_1 di_clk_1 VDD voutn1 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=2*Cu
x11 VSS Vref VSS di_D2_1 di_clk_1 VDD voutn1 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=4*Cu
x12 VSS Vref VSS di_D3_1 di_clk_1 VDD voutn1 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=8*Cu
C1 vinn voutp2 C2 m=1
C2 vinp voutn2 C2 m=1
C1c net2 voutp2 Cucomp m=1
C1d net4 voutn2 Cucomp m=1
x14 VDD di_clk_2 VSS voutp2 Vcm clk_2_n transmission_gate_lv_wo_dummy W_P=1.0u L_P=0.13u W_N=1.0u L_N=0.13u
x15 VDD di_clk_2 VSS voutn2 Vcm clk_2_n transmission_gate_lv_wo_dummy W_P=1.0u L_P=0.13u W_N=1.0u L_N=0.13u
x17 Vref VSS VSS di_D1_2 di_clk_2 VDD voutp2 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=2*Cu
x18 Vref VSS VSS di_D2_2 di_clk_2 VDD voutp2 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=4*Cu
x16 Vref VSS VSS di_D0_2 di_clk_2 VDD voutp2 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=Cu
x19 Vref VSS VSS di_D3_2 di_clk_2 VDD voutp2 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=8*Cu
x21 VSS Vref VSS di_D0_2 di_clk_2 VDD voutn2 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=Cu
x22 VSS Vref VSS di_D1_2 di_clk_2 VDD voutn2 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=2*Cu
x23 VSS Vref VSS di_D2_2 di_clk_2 VDD voutn2 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=4*Cu
x24 VSS Vref VSS di_D3_2 di_clk_2 VDD voutn2 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=8*Cu
x8 VDD di_clk_1 VSS net3 VSS Vref spdt_switch W_P_TG=W_P_SPDT L_P_TG=L_P_SPDT W_N_TG=W_N_SPDT L_N_TG=L_N_SPDT
x13 VDD di_clk_1 VSS net1 Vref VSS spdt_switch W_P_TG=W_P_SPDT L_P_TG=L_P_SPDT W_N_TG=W_N_SPDT L_N_TG=L_N_SPDT
x20 VDD di_clk_2 VSS net2 VSS Vref spdt_switch W_P_TG=W_P_SPDT L_P_TG=L_P_SPDT W_N_TG=W_N_SPDT L_N_TG=L_N_SPDT
x25 VDD di_clk_2 VSS net4 Vref VSS spdt_switch W_P_TG=W_P_SPDT L_P_TG=L_P_SPDT W_N_TG=W_N_SPDT L_N_TG=L_N_SPDT
x26 VDD di_clk_2 clk_2_n VSS inverter_lv W_P=W_P_SPDT L_P=L_P_SPDT W_N=W_N_SPDT L_N=L_N_SPDT
.ends


* expanding   symbol:  top_level/auxiliary/input_hardware.sym # of pins=23
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/top_level/auxiliary/input_hardware.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/top_level/auxiliary/input_hardware.sch
.subckt input_hardware VDD_IO di_clock di_control_mode do_clock do_control_mode VSS di_reset_n do_reset_n di_signal_select_in
+ do_signal_select_in do_enable do_trigger_start_sampling di_trigger_start_sampling di_enable do_select_tbs_delta_steps di_select_tbs_delta_steps
+ do_trigger_start_mode di_trigger_start_mode di_adaptive_mode do_uart_rx do_adaptive_mode di_uart_rx VDD_DIG
*.ipin di_clock
*.ipin di_reset_n
*.ipin di_uart_rx
*.ipin di_trigger_start_sampling
*.ipin di_trigger_start_mode
*.ipin di_adaptive_mode
*.ipin di_control_mode
*.ipin di_signal_select_in
*.ipin di_enable
*.ipin di_select_tbs_delta_steps
*.opin do_clock
*.iopin VDD_IO
*.iopin VDD_DIG
*.opin do_trigger_start_sampling
*.opin do_control_mode
*.opin do_enable
*.opin do_reset_n
*.opin do_trigger_start_mode
*.opin do_adaptive_mode
*.opin do_signal_select_in
*.opin do_select_tbs_delta_steps
*.opin do_uart_rx
*.iopin VSS
x6 VDD_IO net2 di_clock VSS schmitt_trigger W_P_ST=3.0u L_P_ST=0.50u W_N_ST=1.0u L_N_ST=0.50u R=4
x7 VDD_DIG net2 do_clock VSS VDD_IO level_down_shifter W_P_HV=3.0u L_P_HV=0.50u W_N_HV=1.0u L_N_HV=0.50u W_P_LV=3.0u L_P_LV=0.13u
+ W_N_LV=10.0u L_N_LV=0.13u
x10 VDD_IO net3 di_reset_n VSS schmitt_trigger W_P_ST=3.0u L_P_ST=0.50u W_N_ST=1.0u L_N_ST=0.50u R=4
x11 VDD_DIG net3 do_reset_n VSS VDD_IO level_down_shifter W_P_HV=3.0u L_P_HV=0.50u W_N_HV=1.0u L_N_HV=0.50u W_P_LV=3.0u
+ L_P_LV=0.13u W_N_LV=10.0u L_N_LV=0.13u
x12 VDD_IO net4 di_trigger_start_sampling VSS schmitt_trigger W_P_ST=3.0u L_P_ST=0.50u W_N_ST=1.0u L_N_ST=0.50u R=4
x13 VDD_DIG net4 do_trigger_start_sampling VSS VDD_IO level_down_shifter W_P_HV=3.0u L_P_HV=0.50u W_N_HV=1.0u L_N_HV=0.50u
+ W_P_LV=3.0u L_P_LV=0.13u W_N_LV=10.0u L_N_LV=0.13u
x14 VDD_IO net5 di_trigger_start_mode VSS schmitt_trigger W_P_ST=3.0u L_P_ST=0.50u W_N_ST=1.0u L_N_ST=0.50u R=4
x15 VDD_DIG net5 do_trigger_start_mode VSS VDD_IO level_down_shifter W_P_HV=3.0u L_P_HV=0.50u W_N_HV=1.0u L_N_HV=0.50u W_P_LV=3.0u
+ L_P_LV=0.13u W_N_LV=10.0u L_N_LV=0.13u
x16 VDD_IO net1 di_adaptive_mode VSS schmitt_trigger W_P_ST=3.0u L_P_ST=0.50u W_N_ST=1.0u L_N_ST=0.50u R=4
x17 VDD_DIG net1 do_adaptive_mode VSS VDD_IO level_down_shifter W_P_HV=3.0u L_P_HV=0.50u W_N_HV=1.0u L_N_HV=0.50u W_P_LV=3.0u
+ L_P_LV=0.13u W_N_LV=10.0u L_N_LV=0.13u
x18 VDD_IO net6 di_control_mode VSS schmitt_trigger W_P_ST=3.0u L_P_ST=0.50u W_N_ST=1.0u L_N_ST=0.50u R=4
x19 VDD_DIG net6 do_control_mode VSS VDD_IO level_down_shifter W_P_HV=3.0u L_P_HV=0.50u W_N_HV=1.0u L_N_HV=0.50u W_P_LV=3.0u
+ L_P_LV=0.13u W_N_LV=10.0u L_N_LV=0.13u
x20 VDD_IO net7 di_signal_select_in VSS schmitt_trigger W_P_ST=3.0u L_P_ST=0.50u W_N_ST=1.0u L_N_ST=0.50u R=4
x21 VDD_DIG net7 do_signal_select_in VSS VDD_IO level_down_shifter W_P_HV=3.0u L_P_HV=0.50u W_N_HV=1.0u L_N_HV=0.50u W_P_LV=3.0u
+ L_P_LV=0.13u W_N_LV=10.0u L_N_LV=0.13u
x22 VDD_IO net8 di_enable VSS schmitt_trigger W_P_ST=3.0u L_P_ST=0.50u W_N_ST=1.0u L_N_ST=0.50u R=4
x23 VDD_DIG net8 do_enable VSS VDD_IO level_down_shifter W_P_HV=3.0u L_P_HV=0.50u W_N_HV=1.0u L_N_HV=0.50u W_P_LV=3.0u
+ L_P_LV=0.13u W_N_LV=10.0u L_N_LV=0.13u
x24 VDD_IO net9 di_select_tbs_delta_steps VSS schmitt_trigger W_P_ST=3.0u L_P_ST=0.50u W_N_ST=1.0u L_N_ST=0.50u R=4
x25 VDD_DIG net9 do_select_tbs_delta_steps VSS VDD_IO level_down_shifter W_P_HV=3.0u L_P_HV=0.50u W_N_HV=1.0u L_N_HV=0.50u
+ W_P_LV=3.0u L_P_LV=0.13u W_N_LV=10.0u L_N_LV=0.13u
x26 VDD_IO net10 di_uart_rx VSS schmitt_trigger W_P_ST=3.0u L_P_ST=0.50u W_N_ST=1.0u L_N_ST=0.50u R=4
x27 VDD_DIG net10 do_uart_rx VSS VDD_IO level_down_shifter W_P_HV=3.0u L_P_HV=0.50u W_N_HV=1.0u L_N_HV=0.50u W_P_LV=3.0u
+ L_P_LV=0.13u W_N_LV=10.0u L_N_LV=0.13u
.ends


* expanding   symbol:  top_level/auxiliary/output_hardware.sym # of pins=11
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/top_level/auxiliary/output_hardware.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/top_level/auxiliary/output_hardware.sch
.subckt output_hardware di_uart_tx do_uart_tx do_idle_led di_idle_led do_overflow_led di_overflow_led di_underflow_led
+ do_underflow_led VDD_IO VSS VDD_DIG
*.opin do_uart_tx
*.opin do_idle_led
*.opin do_overflow_led
*.opin do_underflow_led
*.iopin VSS
*.iopin VDD_IO
*.iopin VDD_DIG
*.ipin di_idle_led
*.ipin di_overflow_led
*.ipin di_underflow_led
*.ipin di_uart_tx
x8 VDD_IO di_uart_tx do_uart_tx VSS VDD_DIG level_up_shifter W_P_HV=3.0u L_P_HV=0.50u W_N_HV=10.0u L_N_HV=0.50u W_P_LV=1.0u
+ L_P_LV=0.13u W_N_LV=1.0u L_N_LV=0.13u
x9 VDD_IO di_idle_led do_idle_led VSS VDD_DIG level_up_shifter W_P_HV=3.0u L_P_HV=0.50u W_N_HV=10.0u L_N_HV=0.50u W_P_LV=1.0u
+ L_P_LV=0.13u W_N_LV=1.0u L_N_LV=0.13u
x28 VDD_IO di_overflow_led do_overflow_led VSS VDD_DIG level_up_shifter W_P_HV=3.0u L_P_HV=0.50u W_N_HV=10.0u L_N_HV=0.50u
+ W_P_LV=1.0u L_P_LV=0.13u W_N_LV=1.0u L_N_LV=0.13u
x29 VDD_IO di_underflow_led do_underflow_led VSS VDD_DIG level_up_shifter W_P_HV=3.0u L_P_HV=0.50u W_N_HV=10.0u L_N_HV=0.50u
+ W_P_LV=1.0u L_P_LV=0.13u W_N_LV=1.0u L_N_LV=0.13u
.ends


* expanding   symbol:  top_level/auxiliary/esd_protection.sym # of pins=4
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/top_level/auxiliary/esd_protection.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/top_level/auxiliary/esd_protection.sch
.subckt esd_protection VDD vin vout VSS
*.iopin VDD
*.iopin VSS
*.ipin vin
*.opin vout
R1 vin vout 10k m=1
XD1 VDD vout VSS diodevdd_4kv m=1
XD2 VDD vout VSS diodevss_4kv m=1
.ends


* expanding   symbol:  top_level/auxiliary/buffers.sym # of pins=50
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/top_level/auxiliary/buffers.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/top_level/auxiliary/buffers.sch
.subckt buffers VDD_DIG di_phi_dac_lower do_phi_bias_1 di_phi_dac_upper di_phi_cmfb_1 do_phi_dac_lower do_phi_cmfb_1 di_phi_bias_1
+ do_phi_dac_upper VSS di_dac_D0_lower do_dac_D0_lower di_phi_cmfb_2 do_phi_bias_2 di_phi_bias_2 di_dac_D0_upper do_dac_D0_upper do_phi_cmfb_2
+ di_dac_D1_upper do_phi_R_1 di_phi_R_1 do_en_cap_1 do_dac_D1_lower do_dac_D1_upper di_dac_D1_lower di_en_cap_1 di_dac_D2_upper do_phi_R_2
+ di_phi_R_2 do_en_cap_2 do_dac_D2_lower di_en_cap_2 di_dac_D2_lower do_dac_D2_upper do_bio_amp_en do_en_cap_3 di_en_cap_3 di_bio_amp_en
+ do_dac_D3_upper do_dac_D3_lower di_dac_D3_lower di_dac_D3_upper di_phi_comp do_phi_vcm_generator_1 di_phi_vcm_generator_1 do_spdt_ctrl
+ di_spdt_ctrl do_phi_comp do_phi_vcm_generator_2 di_phi_vcm_generator_2
*.iopin VDD_DIG
*.iopin VSS
*.ipin di_phi_dac_upper
*.ipin di_dac_D0_upper
*.ipin di_dac_D1_upper
*.ipin di_dac_D2_upper
*.ipin di_dac_D3_upper
*.opin do_phi_dac_upper
*.opin do_dac_D0_upper
*.opin do_dac_D1_upper
*.opin do_dac_D2_upper
*.opin do_dac_D3_upper
*.ipin di_phi_dac_lower
*.ipin di_dac_D0_lower
*.ipin di_dac_D1_lower
*.ipin di_dac_D2_lower
*.ipin di_dac_D3_lower
*.opin do_phi_dac_lower
*.opin do_dac_D0_lower
*.opin do_dac_D1_lower
*.opin do_dac_D2_lower
*.opin do_dac_D3_lower
*.ipin di_phi_vcm_generator_1
*.opin do_phi_vcm_generator_1
*.ipin di_phi_vcm_generator_2
*.opin do_phi_vcm_generator_2
*.ipin di_phi_cmfb_1
*.opin do_phi_cmfb_1
*.ipin di_phi_cmfb_2
*.opin do_phi_cmfb_2
*.ipin di_phi_comp
*.opin do_phi_comp
*.ipin di_phi_bias_1
*.opin do_phi_bias_1
*.ipin di_en_cap_2
*.opin do_en_cap_2
*.ipin di_en_cap_1
*.opin do_en_cap_1
*.ipin di_spdt_ctrl
*.opin do_spdt_ctrl
*.ipin di_phi_bias_2
*.opin do_phi_bias_2
*.ipin di_phi_R_1
*.opin do_phi_R_1
*.ipin di_phi_R_2
*.opin do_phi_R_2
*.ipin di_en_cap_3
*.opin do_en_cap_3
*.ipin di_bio_amp_en
*.opin do_bio_amp_en
x3 VDD_DIG di_dac_D1_upper do_dac_D1_upper VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x4 VDD_DIG di_dac_D2_upper do_dac_D2_upper VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x1 VDD_DIG di_phi_dac_upper do_phi_dac_upper VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x2 VDD_DIG di_dac_D0_upper do_dac_D0_upper VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x5 VDD_DIG di_dac_D3_upper do_dac_D3_upper VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x6 VDD_DIG di_dac_D1_lower do_dac_D1_lower VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x7 VDD_DIG di_dac_D2_lower do_dac_D2_lower VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x8 VDD_DIG di_phi_dac_lower do_phi_dac_lower VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x9 VDD_DIG di_dac_D0_lower do_dac_D0_lower VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x10 VDD_DIG di_dac_D3_lower do_dac_D3_lower VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x11 VDD_DIG di_phi_vcm_generator_1 do_phi_vcm_generator_1 VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x12 VDD_DIG di_phi_vcm_generator_2 do_phi_vcm_generator_2 VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x13 VDD_DIG di_phi_cmfb_1 do_phi_cmfb_1 VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x14 VDD_DIG di_phi_cmfb_2 do_phi_cmfb_2 VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x15 VDD_DIG di_phi_comp do_phi_comp VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x16 VDD_DIG di_phi_bias_1 do_phi_bias_1 VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x17 VDD_DIG di_en_cap_2 do_en_cap_2 VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x18 VDD_DIG di_en_cap_1 do_en_cap_1 VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x19 VDD_DIG di_spdt_ctrl do_spdt_ctrl VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x20 VDD_DIG di_phi_bias_2 do_phi_bias_2 VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x21 VDD_DIG di_phi_R_1 do_phi_R_1 VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x22 VDD_DIG di_phi_R_2 do_phi_R_2 VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x23 VDD_DIG di_en_cap_3 do_en_cap_3 VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
x24 VDD_DIG di_bio_amp_en do_bio_amp_en VSS buffer_lv W_P_INV=1.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
.ends


* expanding   symbol:  bio_amplifier/sc_fb_resistor/sc_fb_resistor.sym # of pins=6
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/bio_amplifier/sc_fb_resistor/sc_fb_resistor.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/bio_amplifier/sc_fb_resistor/sc_fb_resistor.sch
.subckt sc_fb_resistor sc_fb_a sc_fb_b di_phi_2 di_phi_1 VDD VSS  W_P_FB=1.0u L_P_FB=0.13u W_N_FB=1.0u L_N_FB=0.13u Cs=4f
*.iopin VSS
*.iopin VDD
*.iopin sc_fb_a
*.iopin sc_fb_b
*.ipin di_phi_1
*.ipin di_phi_2
x1 VDD di_phi_1 VSS net1 sc_fb_a di_phi_1_n transmission_gate_lv_wo_dummy W_P=W_P_FB L_P=L_P_FB W_N=W_N_FB L_N=L_N_FB
x2 VDD di_phi_2 VSS net2 net1 di_phi_2_n transmission_gate_lv_wo_dummy W_P=W_P_FB L_P=L_P_FB W_N=W_N_FB L_N=L_N_FB
x3 VDD di_phi_1 VSS net3 net2 di_phi_1_n transmission_gate_lv_wo_dummy W_P=W_P_FB L_P=L_P_FB W_N=W_N_FB L_N=L_N_FB
x4 VDD di_phi_2 VSS net4 net3 di_phi_2_n transmission_gate_lv_wo_dummy W_P=W_P_FB L_P=L_P_FB W_N=W_N_FB L_N=L_N_FB
x5 VDD di_phi_1 VSS net5 net4 di_phi_1_n transmission_gate_lv_wo_dummy W_P=W_P_FB L_P=L_P_FB W_N=W_N_FB L_N=L_N_FB
x6 VDD di_phi_2 VSS sc_fb_b net5 di_phi_2_n transmission_gate_lv_wo_dummy W_P=W_P_FB L_P=L_P_FB W_N=W_N_FB L_N=L_N_FB
C1 net1 VSS Cs m=1
C2 net2 VSS Cs m=1
C3 net3 VSS Cs m=1
C4 net4 VSS Cs m=1
C5 net5 VSS Cs m=1
x7 VDD di_phi_1 di_phi_1_n VSS inverter_lv W_P=W_P_FB L_P=L_P_FB W_N=W_N_FB L_N=L_N_FB
x8 VDD di_phi_2 di_phi_2_n VSS inverter_lv W_P=W_P_FB L_P=L_P_FB W_N=W_N_FB L_N=L_N_FB
.ends


* expanding   symbol:  programmable_cap/programmable_cap_x3.sym # of pins=7
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/programmable_cap/programmable_cap_x3.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/programmable_cap/programmable_cap_x3.sch
.subckt programmable_cap_x3 VDD di_en_1 VSS di_en_2 vcap_1 vcap_2 di_en_3  W_P_PC=1.0u L_P_PC=0.13u W_N_PC=1.0u L_N_PC=0.13u
+ C1=33p C2=132p C3=165p
*.iopin vcap_1
*.iopin vcap_2
*.ipin di_en_1
*.ipin di_en_2
*.ipin di_en_3
*.iopin VDD
*.iopin VSS
x6 VDD di_en_3 VSS net2 vcap_1 di_en_3_n transmission_gate_lv_wo_dummy W_P=W_P_PC L_P=L_P_PC W_N=W_N_PC L_N=L_N_PC
x5 VDD di_en_2 VSS net3 vcap_1 di_en_2_n transmission_gate_lv_wo_dummy W_P=W_P_PC L_P=L_P_PC W_N=W_N_PC L_N=L_N_PC
x4 VDD di_en_1 VSS net1 vcap_1 di_en_1_n transmission_gate_lv_wo_dummy W_P=W_P_PC L_P=L_P_PC W_N=W_N_PC L_N=L_N_PC
C3 net2 vcap_2 C3 m=1
C2 net3 vcap_2 C2 m=1
C1 net1 vcap_2 C1 m=1
x1 VDD di_en_1 di_en_1_n VSS inverter_lv W_P=W_P_PC L_P=L_P_PC W_N=W_N_PC L_N=L_N_PC
x2 VDD di_en_2 di_en_2_n VSS inverter_lv W_P=W_P_PC L_P=L_P_PC W_N=W_N_PC L_N=L_N_PC
x3 VDD di_en_3 di_en_3_n VSS inverter_lv W_P=W_P_PC L_P=L_P_PC W_N=W_N_PC L_N=L_N_PC
.ends


* expanding   symbol:  bio_amplifier/amplifier_core/amplifier_core.sym # of pins=12
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/bio_amplifier/amplifier_core/amplifier_core.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/bio_amplifier/amplifier_core/amplifier_core.sch
.subckt amplifier_core di_phi_cmfb_1 di_phi_bias_2 di_phi_bias_1 di_phi_cmfb_2 voutp voutn di_amp_core_en vinn vinp VDD VSS Vcm
*.ipin di_phi_cmfb_1
*.ipin di_phi_cmfb_2
*.ipin di_phi_bias_1
*.ipin di_phi_bias_2
*.iopin VDD
*.ipin di_amp_core_en
*.ipin vinp
*.ipin vinn
*.opin voutp
*.opin voutn
*.ipin Vcm
*.iopin VSS
x1 VDD di_amp_core_en amp_core_en_n VSS inverter_lv W_P=3.0u L_P=0.13u W_N=1.0u L_N=0.13u
x2 di_phi_cmfb_1 di_phi_cmfb_2 Vcm VDD voutp voutn net3 net4 VSS di_amp_core_en amp_core_en_n Vbiasc Vbias push_pull_amplifier
x3 di_phi_cmfb_1 di_phi_cmfb_2 VDD vinn vinp VSS Vcm di_amp_core_en amp_core_en_n Vbiasc Vbias net1 net2 net4 net3 telescopic_ota
Cm1 voutp net1 1.5p m=1
Cm2 voutn net2 1.5p m=1
x4 di_phi_bias_2 di_phi_bias_1 VDD VSS Vbiasc Vbias di_amp_core_en bias_circuit_4
.ends


* expanding   symbol:  transmission_gate/transmission_gate_lv_wo_dummy.sym # of pins=6
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/transmission_gate/transmission_gate_lv_wo_dummy.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/transmission_gate/transmission_gate_lv_wo_dummy.sch
.subckt transmission_gate_lv_wo_dummy VDD di_tg_ctrl VSS v_b v_a di_tg_ctrl_n  W_P=1.0u L_P=0.13u W_N=1.0u L_N=0.13u
*.iopin v_a
*.iopin v_b
*.iopin VDD
*.iopin VSS
*.ipin di_tg_ctrl
*.ipin di_tg_ctrl_n
XM1 v_a di_tg_ctrl v_b VSS sg13_lv_nmos w=W_N l=L_N ng=1 m=1
XM2 v_a di_tg_ctrl_n v_b VDD sg13_lv_pmos w=W_P l=L_P ng=1 m=1
.ends


* expanding   symbol:  inverter/inverter_lv.sym # of pins=4
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/inverter/inverter_lv.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/inverter/inverter_lv.sch
.subckt inverter_lv VDD vin vout VSS  W_P=3.0u L_P=0.13u W_N=1.0u L_N=0.13u
*.ipin vin
*.iopin VDD
*.iopin VSS
*.opin vout
XM1 vout vin VDD VDD sg13_lv_pmos w=W_P l=L_P ng=1 m=1
XM2 vout vin VSS VSS sg13_lv_nmos w=W_N l=L_N ng=1 m=1
.ends


* expanding   symbol:  buffer/buffer_lv.sym # of pins=4
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/buffer/buffer_lv.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/buffer/buffer_lv.sch
.subckt buffer_lv VDD vin vout VSS  W_P_INV=3.0u L_P_INV=0.13u W_N_INV=1.0u L_N_INV=0.13u
*.ipin vin
*.iopin VDD
*.iopin VSS
*.opin vout
x1 VDD vin net1 VSS inverter_lv W_P=W_P_INV L_P=L_P_INV W_N=W_N_INV L_N=L_N_INV
x2 VDD net1 vout VSS inverter_lv W_P=W_P_INV L_P=L_P_INV W_N=W_N_INV L_N=L_N_INV
.ends


* expanding   symbol:  comparator/SR_latch/SR_latch.sym # of pins=6
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/comparator/SR_latch/SR_latch.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/comparator/SR_latch/SR_latch.sch
.subckt SR_latch VDD S Qn VSS Q R  W_P_SR=1.0u L_P_SR=0.13u W_N_SR=1.0u L_N_SR=0.13u
*.iopin VDD
*.opin Q
*.iopin VSS
*.ipin S
*.ipin R
*.opin Qn
x1 VDD Q R Qn VSS NOR_gate W_P=W_P_SR L_P=L_P_SR W_N=W_N_SR L_N=L_N_SR
x2 VDD Qn Q S VSS NOR_gate W_P=W_P_SR L_P=L_P_SR W_N=W_N_SR L_N=L_N_SR
.ends


* expanding   symbol:  comparator/discrete_time/Dynamic-biasing/dynamic_biasing_comparator.sym # of pins=8
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/comparator/discrete_time/Dynamic-biasing/dynamic_biasing_comparator.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/comparator/discrete_time/Dynamic-biasing/dynamic_biasing_comparator.sch
.subckt dynamic_biasing_comparator di_clk_n di_clk VDD voutp vinp VSS voutn vinn
*.iopin VDD
*.opin voutp
*.opin voutn
*.ipin di_clk_n
*.iopin VSS
*.ipin vinp
*.ipin vinn
*.ipin di_clk
XM3a vs di_clk vctail VSS sg13_lv_nmos w=1.0u l=0.13u ng=1 m=1
XM12 voutp di_clk_n VSS VSS sg13_lv_nmos w=1.0u l=0.13u ng=1 m=1
XM8 net1 voutn VDD VDD sg13_lv_pmos w=2.0u l=0.13u ng=2 m=1
XM10 voutp voutn VSS VSS sg13_lv_nmos w=1.0u l=0.13u ng=1 m=1
XM11 voutn voutp VSS VSS sg13_lv_nmos w=1.0u l=0.13u ng=1 m=1
XM13 voutn di_clk_n VSS VSS sg13_lv_nmos w=1.0u l=0.13u ng=1 m=1
CPn vcpn VSS 300f m=1
CPp vcpp VSS 300f m=1
XM9 net2 voutp VDD VDD sg13_lv_pmos w=2.0u l=0.13u ng=2 m=1
XM6 voutp vcpn net1 VDD sg13_lv_pmos w=2.0u l=0.13u ng=2 m=1
XM7 voutn vcpp net2 VDD sg13_lv_pmos w=2.0u l=0.13u ng=2 m=1
CTAIL vctail VSS 600f m=1
XM3b vctail di_clk_n VSS VSS sg13_lv_nmos w=1.0u l=0.13u ng=1 m=1
XM1 vcpn vinp vs VSS sg13_lv_nmos w=1.0u l=0.13u ng=1 m=1
XM2 vcpp vinn vs VSS sg13_lv_nmos w=1.0u l=0.13u ng=1 m=1
XM4 vcpn di_clk VDD VDD sg13_lv_pmos w=1.0u l=0.13u ng=1 m=1
XM5 vcpp di_clk VDD VDD sg13_lv_pmos w=1.0u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  dac/unit_cell.sym # of pins=7
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/dac/unit_cell.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/dac/unit_cell.sch
.subckt unit_cell v1 v0 VSS di_cell_en di_clk VDD vtop  W_P_SPDT=1.0u L_P_SPDT=0.13u W_N_SPDT=1.0u L_N_SPDT=0.13u Cu=8f
*.iopin VSS
*.iopin A
*.iopin VDD
*.ipin D
*.iopin B
*.iopin vtop
x1 VDD D VSS net1 A B dac_switch W_P_TG=3.0u L_P_TG=0.13u W_N_TG=1.0u L_N_TG=0.13u
XC1 net1 vtop cap_cmim w=7.0e-6 l=7.0e-6 m=1
.ends


* expanding   symbol:  schmitt_trigger/schmitt_trigger.sym # of pins=4
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/schmitt_trigger/schmitt_trigger.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/schmitt_trigger/schmitt_trigger.sch
.subckt schmitt_trigger VDD vout vin VSS  W_P_ST=3.0u L_P_ST=0.50u W_N_ST=1.0u L_N_ST=0.50u R=4
*.iopin VDD
*.opin vout
*.iopin VSS
*.ipin vin
x1 VDD net2 vout VSS inverter_hv W_P=W_P_ST L_P=L_P_ST W_N=W_N_ST L_N=L_N_ST
XM5 net3 vin VDD VDD sg13_hv_pmos w=W_P_ST l=L_P_ST ng=1 m=1
XM4 net2 vin net3 VDD sg13_hv_pmos w=W_P_ST l=L_P_ST ng=1 m=1
XM6 VSS net2 net3 VDD sg13_hv_pmos w=R*W_P_ST l=L_P_ST ng=1 m=1
XM1 net1 vin VSS VSS sg13_hv_nmos w=W_N_ST l=L_N_ST ng=1 m=1
XM2 net2 vin net1 VSS sg13_hv_nmos w=W_N_ST l=L_N_ST ng=1 m=1
XM3 VDD net2 net1 VSS sg13_hv_nmos w=R*W_N_ST l=L_N_ST ng=1 m=1
.ends


* expanding   symbol:  level_shifter/level_down_shifter.sym # of pins=5
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/level_shifter/level_down_shifter.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/level_shifter/level_down_shifter.sch
.subckt level_down_shifter VDD2 A B VSS VDD1  W_P_HV=3.0u L_P_HV=0.50u W_N_HV=1.0u L_N_HV=0.50u W_P_LV=3.0u L_P_LV=0.13u
+ W_N_LV=10.0u L_N_LV=0.13u
*.ipin A
*.iopin VDD1
*.iopin VSS
*.opin B
*.iopin VDD2
x3 VDD2 T B VSS inverter_lv W_P=W_P_LV L_P=L_P_LV W_N=0.1*W_N_LV L_N=L_N_LV
x1 VDD1 A A! VSS inverter_hv W_P=W_P_HV L_P=L_P_HV W_N=W_N_HV L_N=L_N_HV
x2 VDD1 A! net2 VSS inverter_hv W_P=W_P_HV L_P=L_P_HV W_N=W_N_HV L_N=L_N_HV
XM1 net1 A! VSS VSS sg13_lv_nmos w=W_N_LV l=L_N_LV ng=1 m=1
XM3 net1 T VDD2 VDD2 sg13_lv_pmos w=W_P_LV l=L_P_LV ng=1 m=1
XM2 T net2 VSS VSS sg13_lv_nmos w=W_N_LV l=L_N_LV ng=1 m=1
XM4 T net1 VDD2 VDD2 sg13_lv_pmos w=W_P_LV l=L_P_LV ng=1 m=1
.ends


* expanding   symbol:  level_shifter/level_up_shifter.sym # of pins=5
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/level_shifter/level_up_shifter.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/level_shifter/level_up_shifter.sch
.subckt level_up_shifter VDD2 A B VSS VDD1  W_P_HV=3.0u L_P_HV=0.50u W_N_HV=10.0u L_N_HV=0.50u W_P_LV=1.0u L_P_LV=0.13u
+ W_N_LV=1.0u L_N_LV=0.13u
*.ipin A
*.iopin VDD1
*.iopin VSS
*.opin B
*.iopin VDD2
x1 VDD1 A A! VSS inverter_lv W_P=W_P_LV L_P=L_P_LV W_N=W_N_LV L_N=L_N_LV
XM1 net1 A! VSS VSS sg13_hv_nmos w=W_N_HV l=L_N_HV ng=1 m=1
XM4 T net1 VDD2 VDD2 sg13_hv_pmos w=W_P_HV l=L_P_HV ng=1 m=1
x2 VDD1 A! net2 VSS inverter_lv W_P=W_P_LV L_P=L_P_LV W_N=W_N_LV L_N=L_N_LV
XM3 net1 T VDD2 VDD2 sg13_hv_pmos w=W_P_HV l=L_P_HV ng=1 m=1
XM2 T net2 VSS VSS sg13_hv_nmos w=W_N_HV l=L_N_HV ng=1 m=1
x3 VDD2 T B VSS inverter_hv W_P=W_P_HV L_P=L_P_HV W_N=0.1*W_N_HV L_N=L_N_HV
.ends


* expanding   symbol:  bio_amplifier/amplifier_core/push_pull_amplifier/push_pull_amplifier.sym # of pins=13
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/bio_amplifier/amplifier_core/push_pull_amplifier/push_pull_amplifier.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/bio_amplifier/amplifier_core/push_pull_amplifier/push_pull_amplifier.sch
.subckt push_pull_amplifier di_phi_1 di_phi_2 Vcm VDD voutp voutn vinn vinp VSS di_pp_en di_pp_en_n Vbiasc Vbias
*.ipin vinp
*.ipin vinn
*.opin voutp
*.opin voutn
*.iopin VDD
*.iopin VSS
*.ipin di_phi_1
*.ipin di_phi_2
*.ipin Vcm
*.ipin di_pp_en
*.ipin di_pp_en_n
*.ipin Vbias
*.ipin Vbiasc
xM12 voutn Vb VDD VDD sg13g2_lv_pmos_stacked_x4 W_P=4.0u L_P=40.0u NG_P=8 M_P=1
xM10 voutn vinp VSS VSS sg13g2_lv_nmos_stacked_x4 W_N=2.0u L_N=40.0u NG_N=4 M_N=1
xM13 voutp Vb VDD VDD sg13g2_lv_pmos_stacked_x4 W_P=4.0u L_P=40.0u NG_P=8 M_P=1
xM11 voutp vinn VSS VSS sg13g2_lv_nmos_stacked_x4 W_N=2.0u L_N=40.0u NG_N=4 M_N=1
xM16 voutn net1 VDD VDD sg13g2_lv_pmos_stacked_x4 W_P=3.0u L_P=40.0u NG_P=6 M_P=1
xM17 net1 net1 VDD VDD sg13g2_lv_pmos_stacked_x4 W_P=1.0u L_P=40.0u NG_P=2 M_P=1
xM18 net1 vinn VSS VSS sg13g2_lv_nmos_stacked_x4 W_N=0.5u L_N=40.0u NG_N=1 M_N=1
xM19 voutp net2 VDD VDD sg13g2_lv_pmos_stacked_x4 W_P=3.0u L_P=40.0u NG_P=6 M_P=1
xM20 net2 net2 VDD VDD sg13g2_lv_pmos_stacked_x4 W_P=1.0u L_P=40.0u NG_P=2 M_P=1
xM21 net2 vinp VSS VSS sg13g2_lv_nmos_stacked_x4 W_N=0.5u L_N=40.0u NG_N=1 M_N=1
x1 Vcm net3 di_phi_1 di_phi_2 VDD voutp VSS Vb voutn sc_cmfb_output W_P_CMFB=2.0u L_P_CMFB=0.5u W_N_CMFB=2.0u L_N_CMFB=0.5u
+ W_P_CMFB_D=1.0u W_N_CMFB_D=1.0u C1=100f a=9
xM15 net4 net3 VDD VDD sg13g2_lv_pmos_stacked_x4 W_P=2.0u L_P=40.0u NG_P=4 M_P=1
Vmeas3 net4 net5 0
.save i(vmeas3)
XMpd2 net4 di_pp_en_n net3 VDD sg13_hv_pmos w=1.0u l=0.5u ng=1 m=1
XMpd1 net3 di_pp_en VDD VDD sg13_hv_pmos w=1.0u l=0.5u ng=1 m=1
xM14c net5 Vbiasc VSS net6 sg13g2_lv_nmos_stacked_x2 W_N=11.5u L_N=20.0u NG_N=23 M_N=1
xM14 net6 Vbias VSS VSS sg13g2_lv_nmos_stacked_x2 W_N=11.5u L_N=20.0u NG_N=23 M_N=1
.ends


* expanding   symbol:  bio_amplifier/amplifier_core/telescopic_ota/telescopic_ota.sym # of pins=15
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/bio_amplifier/amplifier_core/telescopic_ota/telescopic_ota.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/bio_amplifier/amplifier_core/telescopic_ota/telescopic_ota.sch
.subckt telescopic_ota di_phi_1 di_phi_2 VDD vinn vinp VSS Vcm di_tele_en di_tele_en_n Vbiasc Vbias vmiln vmilp voutp voutn
*.ipin di_phi_1
*.ipin di_phi_2
*.ipin vinp
*.ipin vinn
*.opin voutp
*.opin voutn
*.iopin VDD
*.iopin VSS
*.ipin Vcm
*.ipin di_tele_en
*.ipin di_tele_en_n
*.ipin vmilp
*.ipin vmiln
*.ipin Vbias
*.ipin Vbiasc
x1 di_phi_1 di_phi_2 VDD voutp VSS net7 voutn sc_cmfb_input W_P_CMFB=2.0u L_P_CMFB=0.5u W_N_CMFB=2.0u L_N_CMFB=0.5u C1=100f a=9
xM6 net2 Vgs_m56 VDD VDD sg13g2_lv_pmos_stacked_x2 W_P=1.0u L_P=20.0u NG_P=1 M_P=1
xM5 net1 Vgs_m56 VDD VDD sg13g2_lv_pmos_stacked_x2 W_P=8.0u L_P=20.0u NG_P=8 M_P=1
xM5c Vtail net10 net1 net1 sg13g2_lv_pmos_stacked_x2 W_P=8.0u L_P=20.0u NG_P=8 M_P=1
xM7 net6 net6 net5 net5 sg13g2_lv_pmos_stacked_x2 W_P=0.5u L_P=20.0u NG_P=1 M_P=1
XM1 vmiln vinp net3 net5 sg13_lv_pmos w=250.0u l=10.0u ng=250 m=1
XM1c voutn net6 vmiln vmiln sg13_lv_pmos w=15.0u l=10.0u ng=15 m=1
XM2c voutp net6 vmilp vmilp sg13_lv_pmos w=15.0u l=10.0u ng=15 m=1
XM2 vmilp vinn net4 net5 sg13_lv_pmos w=250.0u l=10.0u ng=250 m=1
xM3 voutn net7 VSS VSS sg13g2_lv_nmos_stacked_x4 W_N=1.5u L_N=40.0u NG_N=1 M_N=1
xM4 voutp net7 VSS VSS sg13g2_lv_nmos_stacked_x4 W_N=1.5u L_N=40.0u NG_N=1 M_N=1
Vmeas net9 net3 0
.save i(vmeas)
Vmeas1 net9 net4 0
.save i(vmeas1)
Vmeas2 net9 net5 0
.save i(vmeas2)
xM6c net8 net10 net2 net2 sg13g2_lv_pmos_stacked_x2 W_P=1.0u L_P=20.0u NG_P=1 M_P=1
XMpd4 Vcm di_tele_en_n net10 VDD sg13_hv_pmos w=1.0u l=0.5u ng=1 m=1
XMdec1 VDD Vgs_m56 VDD VDD sg13_lv_pmos w=10.0u l=40.0u ng=10 m=1
XMpd3 net10 di_tele_en VDD VDD sg13_hv_pmos w=1.0u l=0.5u ng=1 m=1
XMpd2 net8 di_tele_en_n Vgs_m56 VDD sg13_hv_pmos w=1.0u l=0.5u ng=1 m=1
XMpd1 Vgs_m56 di_tele_en VDD VDD sg13_hv_pmos w=1.0u l=0.5u ng=1 m=1
XMdec3 VDD net10 VDD VDD sg13_lv_pmos w=10.0u l=40.0u ng=10 m=1
Vmeas3 net8 net12 0
.save i(vmeas3)
Vmeas4 net6 net14 0
.save i(vmeas4)
xM8c net12 Vbiasc VSS net11 sg13g2_lv_nmos_stacked_x2 W_N=20.0u L_N=20.0u NG_N=20 M_N=1
xM8 net11 Vbias VSS VSS sg13g2_lv_nmos_stacked_x2 W_N=20.0u L_N=20.0u NG_N=20 M_N=1
xM9c net14 Vbiasc VSS net13 sg13g2_lv_nmos_stacked_x2 W_N=10.0u L_N=20.0u NG_N=10 M_N=1
xM9 net13 Vbias VSS VSS sg13g2_lv_nmos_stacked_x2 W_N=10.0u L_N=20.0u NG_N=10 M_N=1
Vmeas5 Vtail net9 0
.save i(vmeas5)
.ends


* expanding   symbol:  bio_amplifier/amplifier_core/bias_circuit/bias_circuit_4/bias_circuit_4.sym # of pins=7
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/bio_amplifier/amplifier_core/bias_circuit/bias_circuit_4/bias_circuit_4.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/bio_amplifier/amplifier_core/bias_circuit/bias_circuit_4/bias_circuit_4.sch
.subckt bias_circuit_4 di_phi_2 di_phi_1 VDD VSS Vbiasc Vbias di_bias_en
*.ipin di_phi_1
*.ipin di_phi_2
*.iopin VDD
*.iopin VSS
*.opin Vbias
*.ipin di_bias_en
*.opin Vbiasc
x2 Vres VSS di_phi_2 di_phi_1 VDD VSS sc_bias_resistor W_P_R=1.0u L_P_R=0.13u W_N_R=1.0u L_N_R=0.13u Cs=1.8p
XMDEC1 net1 Vbias net1 net1 sg13_lv_nmos w=100.0u l=40.0u ng=100 m=1
VIref net3 net5 0
.save i(viref)
VIout net6 Vbiasc 0
.save i(viout)
x1 VDD di_bias_en bias_en_n VSS inverter_lv W_P=1.0u L_P=0.13u W_N=1.0u L_N=0.13u
XMPD1 Vgs_m34 di_bias_en net2 net2 sg13_lv_pmos w=1.0u l=0.13u ng=1 m=1
XMPD2 net3 bias_en_n Vgs_m34 net2 sg13_lv_pmos w=1.0u l=0.13u ng=1 m=1
VIref5 net1 VSS 0
.save i(viref5)
VIdd VDD net2 0
.save i(vidd)
xM1 net4 Vbias VSS Vres sg13g2_lv_nmos_stacked_x2 W_N=20.0u L_N=20.0u NG_N=20 M_N=1
xM1c net5 Vbiasc VSS net4 sg13g2_lv_nmos_stacked_x2 W_N=5.0u L_N=20.0u NG_N=5 M_N=1
xM2 Vbias Vbias VSS VSS sg13g2_lv_nmos_stacked_x2 W_N=5.0u L_N=20.0u NG_N=5 M_N=1
xM2c Vbiasc Vbiasc VSS Vbias sg13g2_lv_nmos_stacked_x2 W_N=5.0u L_N=20.0u NG_N=5 M_N=1
XMDEC2 net2 Vgs_m34 net2 net2 sg13_lv_pmos w=25.0u l=40.0u ng=25 m=1
xM3 net3 Vgs_m34 net2 net2 sg13g2_lv_pmos_stacked_x4 W_P=20.0u L_P=40.0u NG_P=20 M_P=1
xM4 net6 Vgs_m34 net2 net2 sg13g2_lv_pmos_stacked_x4 W_P=20.0u L_P=40.0u NG_P=20 M_P=1
XMDEC3 VSS Vres VSS VSS sg13_lv_nmos w=43.0u l=40.0u ng=43 m=1
xMSU2 Vsu net8 VSS VSS sg13g2_lv_nmos_stacked_x4 W_N=1.0u L_N=40.0u NG_N=1 M_N=1
xMSU1 net7 Vsu VSS net8 sg13g2_lv_nmos_stacked_x4 W_N=1.0u L_N=40.0u NG_N=1 M_N=1
Vmeas1 net3 net7 0
.save i(vmeas1)
Vmeas2 Vbias net8 0
.save i(vmeas2)
CSU1 net9 Vsu 35f m=1
XMPD6 Vsu di_bias_en net9 net9 sg13_lv_pmos w=1.0u l=0.13u ng=1 m=1
XMPD7 Vsu bias_en_n VSS VSS sg13_lv_nmos w=1.0u l=0.13u ng=1 m=1
XMPD5 net9 bias_en_n net2 net2 sg13_lv_pmos w=1.0u l=0.13u ng=1 m=1
XMPD3 Vbias bias_en_n VSS VSS sg13_lv_nmos w=1.0u l=0.13u ng=1 m=1
XMPD4 Vbias bias_en_n VSS VSS sg13_lv_nmos w=1.0u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  comparator/NOR_gate/NOR_gate.sym # of pins=5
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/comparator/NOR_gate/NOR_gate.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/comparator/NOR_gate/NOR_gate.sch
.subckt NOR_gate VDD C A B VSS  W_P=1.0u L_P=0.13u W_N=0.5u L_N=0.13u
*.iopin VDD
*.opin C
*.iopin VSS
*.ipin A
*.ipin B
XM1 C A VSS VSS sg13_lv_nmos w=W_N l=L_N ng=1 m=1
XM2 C B VSS VSS sg13_lv_nmos w=W_N l=L_N ng=1 m=1
XM3 C B net1 VDD sg13_lv_pmos w=W_P l=L_P ng=1 m=1
XM4 net1 A VDD VDD sg13_lv_pmos w=W_P l=L_P ng=1 m=1
XM5 C A net2 VDD sg13_lv_pmos w=W_P l=L_P ng=1 m=1
XM6 net2 B VDD VDD sg13_lv_pmos w=W_P l=L_P ng=1 m=1
.ends


* expanding   symbol:  dac_icms_cell/dac_switch.sym # of pins=6
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/dac_icms_cell/dac_switch.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/dac_icms_cell/dac_switch.sch
.subckt dac_switch VDD di_spdt_ctrl VSS v_c v_b v_a  W_P_TG=3.0u L_P_TG=0.13u W_N_TG=1.0u L_N_TG=0.13u
*.iopin v_a
*.iopin v_c
*.iopin VDD
*.iopin VSS
*.ipin di_spdt_ctrl
*.iopin v_b
x1 VDD di_spdt_ctrl VSS v_c v_a di_spdt_ctrl_n transmission_gate_lv_wo_dummy W_P=W_P_TG L_P=L_P_TG W_N=W_N_TG L_N=L_N_TG
x8 VDD di_spdt_ctrl di_spdt_ctrl_n VSS inverter_lv W_P=W_P_TG L_P=L_P_TG W_N=W_N_TG L_N=L_N_TG
XM5 net2 di_spdt_ctrl_n VSS VSS sg13_hv_nmos w=0.3u l=0.6u ng=1 m=1
XM4 net1 di_spdt_ctrl VDD VDD sg13_hv_pmos w=0.3u l=0.6u ng=1 m=1
XM1 v_c v_b net2 VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM3 v_c v_b net1 VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  inverter/inverter_hv.sym # of pins=4
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/inverter/inverter_hv.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/inverter/inverter_hv.sch
.subckt inverter_hv VDD vin vout VSS  W_P=3.0u L_P=0.50u W_N=1.0u L_N=0.50u
*.ipin vin
*.iopin VDD
*.iopin VSS
*.opin vout
XM1 vout vin VDD VDD sg13_hv_pmos w=W_P l=L_P ng=1 m=1
XM2 vout vin VSS VSS sg13_hv_nmos w=W_N l=L_N ng=1 m=1
.ends


* expanding   symbol:  stacked_transistors/sg13g2_lv_pmos_stacked/sg13g2_lv_pmos_stacked_x4.sym # of pins=4
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/stacked_transistors/sg13g2_lv_pmos_stacked/sg13g2_lv_pmos_stacked_x4.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/stacked_transistors/sg13g2_lv_pmos_stacked/sg13g2_lv_pmos_stacked_x4.sch
.subckt sg13g2_lv_pmos_stacked_x4 D G B S  W_P=1.0u L_P=0.45u NG_P=1 M_P=1
*.iopin D
*.iopin S
*.iopin G
*.iopin B
XM1 net1 G S B sg13_lv_pmos w=W_P l=L_P/4 ng=NG_P m=M_P
XM2 net3 G net1 B sg13_lv_pmos w=W_P l=L_P/4 ng=NG_P m=M_P
XM3 net2 G net3 B sg13_lv_pmos w=W_P l=L_P/4 ng=NG_P m=M_P
XM4 D G net2 B sg13_lv_pmos w=W_P l=L_P/4 ng=NG_P m=M_P
.ends


* expanding   symbol:  stacked_transistors/sg13g2_lv_nmos_stacked/sg13g2_lv_nmos_stacked_x4.sym # of pins=4
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/stacked_transistors/sg13g2_lv_nmos_stacked/sg13g2_lv_nmos_stacked_x4.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/stacked_transistors/sg13g2_lv_nmos_stacked/sg13g2_lv_nmos_stacked_x4.sch
.subckt sg13g2_lv_nmos_stacked_x4 D G B S  W_N=1.0u L_N=0.45u NG_N=1 M_N=1
*.iopin D
*.iopin S
*.iopin G
*.iopin B
XM1 net1 G S B sg13_lv_nmos w=W_N l=L_N/4 ng=NG_N m=M_N
XM2 net3 G net1 B sg13_lv_nmos w=W_N l=L_N/4 ng=NG_N m=M_N
XM3 net2 G net3 B sg13_lv_nmos w=W_N l=L_N/4 ng=NG_N m=M_N
XM4 D G net2 B sg13_lv_nmos w=W_N l=L_N/4 ng=NG_N m=M_N
.ends


* expanding   symbol:  bio_amplifier/amplifier_core/sc_cmfb/sc_cmfb_output.sym # of pins=9
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/bio_amplifier/amplifier_core/sc_cmfb/sc_cmfb_output.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/bio_amplifier/amplifier_core/sc_cmfb/sc_cmfb_output.sch
.subckt sc_cmfb_output Vcmref Vbias di_phi_1 di_phi_2 VDD Voutp VSS Vb Voutn  W_P_CMFB=2.0u L_P_CMFB=0.5u W_N_CMFB=2.0u
+ L_N_CMFB=0.5u W_P_CMFB_D=1.0u W_N_CMFB_D=1.0u C1=100f a=9
*.iopin VSS
*.iopin VDD
*.iopin Vb
*.iopin Voutp
*.iopin Voutn
*.iopin Vbias
*.iopin Vcmref
*.ipin di_phi_1
*.ipin di_phi_2
x1 VDD di_phi_2 VSS net1 Voutp di_phi_2_n transmission_gate_lv_wo_dummy W_P=W_P_CMFB L_P=L_P_CMFB W_N=W_N_CMFB L_N=L_N_CMFB
C1 Voutp Vb {a*C1} m=1
x2 VDD di_phi_2 VSS net3 Vb di_phi_2_n transmission_gate_lv_wo_dummy W_P=W_P_CMFB L_P=L_P_CMFB W_N=W_N_CMFB L_N=L_N_CMFB
x3 VDD di_phi_2 VSS net2 Voutn di_phi_2_n transmission_gate_lv_wo_dummy W_P=W_P_CMFB L_P=L_P_CMFB W_N=W_N_CMFB L_N=L_N_CMFB
C2 Vb Voutn {a*C1} m=1
C3 net1 net3 C1 m=1
C4 net3 net2 C1 m=1
x7 VDD di_phi_1 di_phi_1_n VSS inverter_lv W_P=W_P_CMFB/2 L_P=L_P_CMFB W_N=W_N_CMFB/2 L_N=L_N_CMFB
x8 VDD di_phi_2 di_phi_2_n VSS inverter_lv W_P=W_P_CMFB/2 L_P=L_P_CMFB W_N=W_N_CMFB/2 L_N=L_N_CMFB
x4 VDD di_phi_1 VSS Vcmref net1 di_phi_1_n transmission_gate_lv_w_dummy W_P=W_P_CMFB L_P=L_P_CMFB W_N=W_N_CMFB L_N=L_N_CMFB
+ W_P_D=W_P_CMFB_D L_P_D=L_P_CMFB W_N_D=W_N_CMFB_D L_N_D=L_N_CMFB
x5 VDD di_phi_1 VSS Vbias net3 di_phi_1_n transmission_gate_lv_w_dummy W_P=W_P_CMFB L_P=L_P_CMFB W_N=W_N_CMFB L_N=L_N_CMFB
+ W_P_D=W_P_CMFB_D L_P_D=L_P_CMFB W_N_D=W_N_CMFB_D L_N_D=L_N_CMFB
x6 VDD di_phi_1 VSS Vcmref net2 di_phi_1_n transmission_gate_lv_w_dummy W_P=W_P_CMFB L_P=L_P_CMFB W_N=W_N_CMFB L_N=L_N_CMFB
+ W_P_D=W_P_CMFB_D L_P_D=L_P_CMFB W_N_D=W_N_CMFB_D L_N_D=L_N_CMFB
.ends


* expanding   symbol:  stacked_transistors/sg13g2_lv_nmos_stacked/sg13g2_lv_nmos_stacked_x2.sym # of pins=4
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/stacked_transistors/sg13g2_lv_nmos_stacked/sg13g2_lv_nmos_stacked_x2.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/stacked_transistors/sg13g2_lv_nmos_stacked/sg13g2_lv_nmos_stacked_x2.sch
.subckt sg13g2_lv_nmos_stacked_x2 D G B S  W_N=1.0u L_N=0.45u NG_N=1 M_N=1
*.iopin D
*.iopin S
*.iopin G
*.iopin B
XM1 net1 G S B sg13_lv_nmos w=W_N l=L_N/2 ng=NG_N m=M_N
XM2 D G net1 B sg13_lv_nmos w=W_N l=L_N/2 ng=NG_N m=M_N
.ends


* expanding   symbol:  bio_amplifier/amplifier_core/sc_cmfb/sc_cmfb_input.sym # of pins=7
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/bio_amplifier/amplifier_core/sc_cmfb/sc_cmfb_input.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/bio_amplifier/amplifier_core/sc_cmfb/sc_cmfb_input.sch
.subckt sc_cmfb_input di_phi_1 di_phi_2 VDD Voutp VSS Vcmfb Voutn  W_P_CMFB=2.0u L_P_CMFB=0.5u W_N_CMFB=2.0u L_N_CMFB=0.5u C1=100f
+ a=9
*.iopin VSS
*.iopin VDD
*.iopin Vcmfb
*.iopin Voutp
*.iopin Voutn
*.ipin di_phi_1
*.ipin di_phi_2
x1 VDD di_phi_2 VSS net1 Voutp di_phi_2_n transmission_gate_lv_wo_dummy W_P=W_P_CMFB L_P=L_P_CMFB W_N=W_N_CMFB L_N=L_N_CMFB
C1 Voutp Vcmfb {a*C1} m=1
x2 VDD di_phi_2 VSS net2 Vcmfb di_phi_2_n transmission_gate_lv_wo_dummy W_P=W_P_CMFB L_P=L_P_CMFB W_N=W_N_CMFB L_N=L_N_CMFB
x3 VDD di_phi_2 VSS net3 Voutn di_phi_2_n transmission_gate_lv_wo_dummy W_P=W_P_CMFB L_P=L_P_CMFB W_N=W_N_CMFB L_N=L_N_CMFB
x4 VDD di_phi_1 VSS net2 net1 di_phi_1_n transmission_gate_lv_wo_dummy W_P=W_P_CMFB L_P=L_P_CMFB W_N=W_N_CMFB L_N=L_N_CMFB
x5 VDD di_phi_1 VSS net2 net3 di_phi_1_n transmission_gate_lv_wo_dummy W_P=W_P_CMFB L_P=L_P_CMFB W_N=W_N_CMFB L_N=L_N_CMFB
C2 Vcmfb Voutn {a*C1} m=1
C3 net1 net2 C1 m=1
C4 net2 net3 C1 m=1
x7 VDD di_phi_1 di_phi_1_n VSS inverter_lv W_P=W_P_CMFB L_P=L_P_CMFB W_N=W_N_CMFB L_N=L_N_CMFB
x6 VDD di_phi_2 di_phi_2_n VSS inverter_lv W_P=W_P_CMFB L_P=L_P_CMFB W_N=W_N_CMFB L_N=L_N_CMFB
.ends


* expanding   symbol:  stacked_transistors/sg13g2_lv_pmos_stacked/sg13g2_lv_pmos_stacked_x2.sym # of pins=4
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/stacked_transistors/sg13g2_lv_pmos_stacked/sg13g2_lv_pmos_stacked_x2.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/stacked_transistors/sg13g2_lv_pmos_stacked/sg13g2_lv_pmos_stacked_x2.sch
.subckt sg13g2_lv_pmos_stacked_x2 D G B S  W_P=1.0u L_P=0.45u NG_P=1 M_P=1
*.iopin D
*.iopin S
*.iopin G
*.iopin B
XM1 net1 G S B sg13_lv_pmos w=W_P l=L_P/2 ng=NG_P m=M_P
XM2 D G net1 B sg13_lv_pmos w=W_P l=L_P/2 ng=NG_P m=M_P
.ends


* expanding   symbol:  bio_amplifier/amplifier_core/bias_circuit/sc_bias_resistor/sc_bias_resistor.sym # of pins=6
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/bio_amplifier/amplifier_core/bias_circuit/sc_bias_resistor/sc_bias_resistor.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/bio_amplifier/amplifier_core/bias_circuit/sc_bias_resistor/sc_bias_resistor.sch
.subckt sc_bias_resistor sc_R_a sc_R_b di_phi_2 di_phi_1 VDD VSS  W_P_R=1.0u L_P_R=0.13u W_N_R=1.0u L_N_R=0.13u Cs=100f
*.iopin VSS
*.iopin VDD
*.iopin sc_R_a
*.iopin sc_R_b
*.ipin di_phi_1
*.ipin di_phi_2
C1 net1 sc_R_b Cs m=1
x1 VDD di_phi_1 VSS net1 sc_R_a di_phi_1_n transmission_gate_lv_wo_dummy W_P=W_P_R L_P=L_P_R W_N=W_N_R L_N=L_N_R
x2 VDD di_phi_2 VSS sc_R_b net1 di_phi_2_n transmission_gate_lv_wo_dummy W_P=W_P_R L_P=L_P_R W_N=W_N_R L_N=L_N_R
C2 net2 sc_R_b Cs m=1
x3 VDD di_phi_2 VSS net2 sc_R_a di_phi_2_n transmission_gate_lv_wo_dummy W_P=W_P_R L_P=L_P_R W_N=W_N_R L_N=L_N_R
x4 VDD di_phi_1 VSS sc_R_b net2 di_phi_1_n transmission_gate_lv_wo_dummy W_P=W_P_R L_P=L_P_R W_N=W_N_R L_N=L_N_R
x5 VDD di_phi_1 di_phi_1_n VSS inverter_lv W_P=W_P_R L_P=L_P_R W_N=W_N_R L_N=L_N_R
x6 VDD di_phi_2 di_phi_2_n VSS inverter_lv W_P=W_P_R L_P=L_P_R W_N=W_N_R L_N=L_N_R
.ends


* expanding   symbol:  transmission_gate/transmission_gate_lv_w_dummy.sym # of pins=6
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/transmission_gate/transmission_gate_lv_w_dummy.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/transmission_gate/transmission_gate_lv_w_dummy.sch
.subckt transmission_gate_lv_w_dummy VDD di_tg_ctrl VSS v_b v_a di_tg_ctrl_n  W_P=2.0u L_P=0.13u W_N=2.0u L_N=0.13u W_P_D=1.0u
+ L_P_D=0.13u W_N_D=1.0u L_N_D=0.13u
*.iopin v_a
*.iopin v_b
*.iopin VDD
*.iopin VSS
*.ipin di_tg_ctrl
*.ipin di_tg_ctrl_n
XM1 v_a di_tg_ctrl v_b VSS sg13_lv_nmos w=W_N l=L_N ng=1 m=1
XM2 v_a di_tg_ctrl_n v_b VDD sg13_lv_pmos w=W_P l=L_P ng=1 m=1
XMdummy2 v_b di_tg_ctrl v_b VDD sg13_lv_pmos w=W_P_D l=L_P_D ng=1 m=1
XMdummy1 v_b di_tg_ctrl_n v_b VSS sg13_lv_nmos w=W_N_D l=L_N_D ng=1 m=1
.ends

.GLOBAL GND
.end
