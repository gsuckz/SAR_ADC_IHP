** sch_path: /foss/designs/SAR_ADC_IHP/xschem/comparator/discrete_time/StrongARM/testbenches/StrongARM_comparator_tb_tran.sch
**.subckt StrongARM_comparator_tb_tran
VDD VDD GND 1.5
V1 clk GND pulse(0 1.5 {tstart} 10p 10p {1/fclk} {1/fphi})
vinn vinn GND {Vcm}
vinp vinp GND {{Vcm} + {delta_vin}}
C1 voutn GND 10f m=1
C2 voutp GND 10f m=1
x1 clk VDD voutp vinp GND voutn vinn StrongARM_comparator
**** begin user architecture code

.lib cornerMOSlv.lib mos_tt
.lib cornerMOShv.lib mos_tt
.lib cornerRES.lib res_typ



.param temp=27
.param fclk=8000000
.param fphi=62500
.param tstart=2n
.param delta_vin = 10m
.param Vcm=0.75
.csparam fclk=fclk
.csparam tstart=tstart
.options savecurrents reltol=1e-3 abstol=1e-12 gmin=1e-15
.control
save all

* Operating Point Analysis
op
remzerovec
write StrongARM_comparator_tb_tran.raw
set appendwrite

* Transient Analysis
* tran 4p 20n
tran 40p 150n
write StrongARM_comparator_tb_tran.raw

* Measure Propagation Delay
* Time from clock rising edge to 90% VDD of voutp
let voutp_limit = 0.9 * 1.5
meas tran tcross WHEN v(voutp)=voutp_limit CROSS=2
let tpd = tcross - tstart
echo Propagation Delay $&tpd s

* Calculate Energy / Conversion
* i_int in As
* energy_conv in Ws = J
let N = 1
let t_conv = 150n
meas tran i_int INTEG i(VDD) from=tstart to=t_conv
let energy_conv = 1.5 * i_int / N

let energy_conv_femto = energy_conv * 1e15
echo Energy / Conversion $&energy_conv_femto fJ/conv

* Plotting
plot v(clk) v(x1.vs) v(voutp) v(voutn)

plot i(VDD)

*quit
.endc

**** end user architecture code
**.ends

* expanding   symbol:  comparator/discrete_time/StrongARM/StrongARM_comparator.sym # of pins=7
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/comparator/discrete_time/StrongARM/StrongARM_comparator.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/comparator/discrete_time/StrongARM/StrongARM_comparator.sch
.subckt StrongARM_comparator di_clk VDD voutp vinp VSS voutn vinn
*.iopin VDD
*.opin voutp
*.iopin VSS
*.opin voutn
*.ipin vinp
*.ipin vinn
*.ipin di_clk
XM1 net1 vinp vs VSS sg13_lv_nmos w=1.0u l=0.13u ng=1 m=1
XM2 net2 vinn vs VSS sg13_lv_nmos w=1.0u l=0.13u ng=1 m=1
XM3 voutn voutp net1 VSS sg13_lv_nmos w=1.0u l=0.13u ng=1 m=1
XM4 voutp voutn net2 VSS sg13_lv_nmos w=1.0u l=0.13u ng=1 m=1
XM5 voutn voutp VDD VDD sg13_lv_pmos w=1.0u l=0.13u ng=1 m=1
XM6 voutp voutn VDD VDD sg13_lv_pmos w=1.0u l=0.13u ng=1 m=1
XM7 vs di_clk VSS VSS sg13_lv_nmos w=1.0u l=0.13u ng=1 m=1
XM8 voutn di_clk VDD VDD sg13_lv_pmos w=1.0u l=0.13u ng=1 m=1
XM9 net1 di_clk VDD VDD sg13_lv_pmos w=1.0u l=0.13u ng=1 m=1
XM10 voutp di_clk VDD VDD sg13_lv_pmos w=1.0u l=0.13u ng=1 m=1
XM11 net2 di_clk VDD VDD sg13_lv_pmos w=1.0u l=0.13u ng=1 m=1
CPn voutn VSS 300f m=1
CPp voutp VSS 300f m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.end
