** sch_path: /foss/designs/SAR_ADC_IHP/xschem/dac/testbenches/dac_tb_tran.sch
**.subckt dac_tb_tran
VDD VDD GND 1.5
Vclk clk GND pulse(0 1.5 0 1p 1p {1/fclk} {1/fphi})
Vcm Vcm GND 0.75
E4 Vcm vinn net1 GND 0.5
E5 vinp Vcm net1 GND 0.5
E6 net1 GND vind GND 1
vsine vind GND sin(0 1.5 512)
VD0 D0 GND {{D0}*1.5}
VD1 D1 GND {{D1}*1.5}
VD2 D2 GND {{D2}*1.5}
VD3 D3 GND {{D3}*1.5}
C1 voutn2 GND {Cl} m=1
C2 voutp2 GND {Cl} m=1
C3 voutn1 GND {Cl} m=1
C4 voutp1 GND {Cl} m=1
x1 VDD vinp voutp1 voutn1 vinn D0 D1 D2 D3 GND VDD Vcm voutp2 voutn2 clk D0 D1 D2 D3 clk dac W_P_SPDT=1.0u L_P_SPDT=0.13u W_N_SPDT=1.0u
+ L_N_SPDT=0.13u C2={C2} Cu={Cu} Cucomp={Cucomp}
**** begin user architecture code

.lib cornerMOSlv.lib mos_tt
.lib cornerMOShv.lib mos_tt
.lib cornerRES.lib res_typ



.param temp=27
.param C2 = 1024f
.param Cu = 8f
.param Cucomp = 8.1f
* Cl = approx. Cin of DT Comparator
.param Cl = 1.2f
.param W_P = 1.0u
.param L_P = 0.13u
.param W_N = 1.0u
.param L_N = 0.13u
.param fclk=8000000
.csparam fclk = fclk
* Ensure that 1/fphi is an exact multiple of 1/fclk.
* Take approx. Tavg for a good result for sine waves.
* fphi=7812.5, fphi=15625, fphi=31250, fphi=62500, fphi=125000
.param fphi=15625
.param D0 = 1
.param D1 = 1
.param D2 = 1
.param D3 = 0
.options savecurrents klu method=gear reltol=1e-3 abstol=1e-12 gmin=1e-15
.control

save all
* save v(VDD) v(Vcm) v(clk) v(D0) v(D1) v(D2) v(D3) v(vind) v(vinp) v(vinn) v(voutp1) v(voutn1) v(voutp2) v(voutn2)

* User Constants
let tstop = 2m
let tstep = 1/fclk

* Transient Analysis
tran $&tstep $&tstop
write dac_tb_tran.raw
set appendwrite

* Plotting
let vin = vinp - vinn
let vout1 = voutp1 - voutn1
let vout2 = voutp2 - voutn2
plot vin
plot vout1 voutp1 voutn1
plot vout2 voutp2 voutn2

* Measurement of start voltages
meas tran vstart1 FIND vout1 at=150n
meas tran vstart2 FIND vout2 at=150n

* Calculate Power Consumption
* i_int in As
* energy in Ws = J
meas tran i_int INTEG i(VDD) from=0p to=tstop
let energy = 1.5 * i_int
let energy_pico = energy * 1e12
echo Energy $&energy_pico pJ
let power = energy / tstop * 1e9
echo Power Consumption $&power nW

.endc


**** end user architecture code
**.ends

* expanding   symbol:  dac/dac.sym # of pins=20
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/dac/dac.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/dac/dac.sch
.subckt dac VDD vinp voutp1 voutn1 vinn di_D0_2 di_D1_2 di_D2_2 di_D3_2 VSS Vref Vcm voutp2 voutn2 di_clk_2 di_D0_1 di_D1_1
+ di_D2_1 di_D3_1 di_clk_1  W_P_SPDT=1.0u L_P_SPDT=0.13u W_N_SPDT=1.0u L_N_SPDT=0.13u C2=1024f Cu=8f Cucomp=8.1f
*.opin voutp1
*.ipin di_D0_1
*.iopin VSS
*.iopin Vref
*.opin voutn1
*.ipin vinp
*.ipin vinn
*.ipin di_D1_1
*.ipin di_D2_1
*.ipin di_D3_1
*.opin voutp2
*.opin voutn2
*.iopin VDD
*.ipin Vcm
*.ipin di_clk_1
*.ipin di_D3_2
*.ipin di_D2_2
*.ipin di_D1_2
*.ipin di_D0_2
*.ipin di_clk_2
C2a vinp voutp1 C2 m=1
C2b vinn voutn1 C2 m=1
C1a net3 voutp1 Cucomp m=1
C1b net1 voutn1 Cucomp m=1
x2 VDD di_clk_1 VSS voutp1 Vcm clk_1_n transmission_gate_lv_wo_dummy W_P=1.0u L_P=0.13u W_N=1.0u L_N=0.13u
x3 VDD di_clk_1 VSS voutn1 Vcm clk_1_n transmission_gate_lv_wo_dummy W_P=1.0u L_P=0.13u W_N=1.0u L_N=0.13u
x1 VDD di_clk_1 clk_1_n VSS inverter_lv W_P=W_P_SPDT L_P=L_P_SPDT W_N=W_N_SPDT L_N=L_N_SPDT
x5 Vref VSS VSS di_D1_1 di_clk_1 VDD voutp1 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=2*Cu
x6 Vref VSS VSS di_D2_1 di_clk_1 VDD voutp1 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=4*Cu
x4 Vref VSS VSS di_D0_1 di_clk_1 VDD voutp1 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=Cu
x7 Vref VSS VSS di_D3_1 di_clk_1 VDD voutp1 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=8*Cu
x9 VSS Vref VSS di_D0_1 di_clk_1 VDD voutn1 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=Cu
x10 VSS Vref VSS di_D1_1 di_clk_1 VDD voutn1 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=2*Cu
x11 VSS Vref VSS di_D2_1 di_clk_1 VDD voutn1 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=4*Cu
x12 VSS Vref VSS di_D3_1 di_clk_1 VDD voutn1 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=8*Cu
C1 vinn voutp2 C2 m=1
C2 vinp voutn2 C2 m=1
C1c net2 voutp2 Cucomp m=1
C1d net4 voutn2 Cucomp m=1
x14 VDD di_clk_2 VSS voutp2 Vcm clk_2_n transmission_gate_lv_wo_dummy W_P=1.0u L_P=0.13u W_N=1.0u L_N=0.13u
x15 VDD di_clk_2 VSS voutn2 Vcm clk_2_n transmission_gate_lv_wo_dummy W_P=1.0u L_P=0.13u W_N=1.0u L_N=0.13u
x17 Vref VSS VSS di_D1_2 di_clk_2 VDD voutp2 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=2*Cu
x18 Vref VSS VSS di_D2_2 di_clk_2 VDD voutp2 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=4*Cu
x16 Vref VSS VSS di_D0_2 di_clk_2 VDD voutp2 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=Cu
x19 Vref VSS VSS di_D3_2 di_clk_2 VDD voutp2 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=8*Cu
x21 VSS Vref VSS di_D0_2 di_clk_2 VDD voutn2 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=Cu
x22 VSS Vref VSS di_D1_2 di_clk_2 VDD voutn2 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=2*Cu
x23 VSS Vref VSS di_D2_2 di_clk_2 VDD voutn2 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=4*Cu
x24 VSS Vref VSS di_D3_2 di_clk_2 VDD voutn2 unit_cell W_P_SPDT=W_P_SPDT L_P_SPDT=L_P_SPDT W_N_SPDT=W_N_SPDT L_N_SPDT=L_N_SPDT
+ Cu=8*Cu
x8 VDD di_clk_1 VSS net3 VSS Vref spdt_switch W_P_TG=W_P_SPDT L_P_TG=L_P_SPDT W_N_TG=W_N_SPDT L_N_TG=L_N_SPDT
x13 VDD di_clk_1 VSS net1 Vref VSS spdt_switch W_P_TG=W_P_SPDT L_P_TG=L_P_SPDT W_N_TG=W_N_SPDT L_N_TG=L_N_SPDT
x20 VDD di_clk_2 VSS net2 VSS Vref spdt_switch W_P_TG=W_P_SPDT L_P_TG=L_P_SPDT W_N_TG=W_N_SPDT L_N_TG=L_N_SPDT
x25 VDD di_clk_2 VSS net4 Vref VSS spdt_switch W_P_TG=W_P_SPDT L_P_TG=L_P_SPDT W_N_TG=W_N_SPDT L_N_TG=L_N_SPDT
x26 VDD di_clk_2 clk_2_n VSS inverter_lv W_P=W_P_SPDT L_P=L_P_SPDT W_N=W_N_SPDT L_N=L_N_SPDT
.ends


* expanding   symbol:  transmission_gate/transmission_gate_lv_wo_dummy.sym # of pins=6
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/transmission_gate/transmission_gate_lv_wo_dummy.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/transmission_gate/transmission_gate_lv_wo_dummy.sch
.subckt transmission_gate_lv_wo_dummy VDD di_tg_ctrl VSS v_b v_a di_tg_ctrl_n  W_P=1.0u L_P=0.13u W_N=1.0u L_N=0.13u
*.iopin v_a
*.iopin v_b
*.iopin VDD
*.iopin VSS
*.ipin di_tg_ctrl
*.ipin di_tg_ctrl_n
XM1 v_a di_tg_ctrl v_b VSS sg13_lv_nmos w=W_N l=L_N ng=1 m=1
XM2 v_a di_tg_ctrl_n v_b VDD sg13_lv_pmos w=W_P l=L_P ng=1 m=1
.ends


* expanding   symbol:  inverter/inverter_lv.sym # of pins=4
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/inverter/inverter_lv.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/inverter/inverter_lv.sch
.subckt inverter_lv VDD vin vout VSS  W_P=3.0u L_P=0.13u W_N=1.0u L_N=0.13u
*.ipin vin
*.iopin VDD
*.iopin VSS
*.opin vout
XM1 vout vin VDD VDD sg13_lv_pmos w=W_P l=L_P ng=1 m=1
XM2 vout vin VSS VSS sg13_lv_nmos w=W_N l=L_N ng=1 m=1
.ends


* expanding   symbol:  dac/unit_cell.sym # of pins=7
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/dac/unit_cell.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/dac/unit_cell.sch
.subckt unit_cell v1 v0 VSS di_cell_en di_clk VDD vtop  W_P_SPDT=1.0u L_P_SPDT=0.13u W_N_SPDT=1.0u L_N_SPDT=0.13u Cu=8f
*.iopin VSS
*.iopin A
*.iopin VDD
*.ipin D
*.iopin B
*.iopin vtop
x1 VDD D VSS net1 A B dac_switch W_P_TG=3.0u L_P_TG=0.13u W_N_TG=1.0u L_N_TG=0.13u
XC1 net1 vtop cap_cmim w=7.0e-6 l=7.0e-6 m=1
.ends


* expanding   symbol:  spdt_switch/spdt_switch.sym # of pins=6
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/spdt_switch/spdt_switch.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/spdt_switch/spdt_switch.sch
.subckt spdt_switch VDD di_spdt_ctrl VSS v_c v_b v_a  W_P_TG=3.0u L_P_TG=0.13u W_N_TG=1.0u L_N_TG=0.13u
*.iopin v_a
*.iopin v_b
*.iopin v_c
*.iopin VDD
*.iopin VSS
*.ipin di_spdt_ctrl
x1 VDD di_spdt_ctrl VSS v_c v_a di_spdt_ctrl_n transmission_gate_lv_wo_dummy W_P=W_P_TG L_P=L_P_TG W_N=W_N_TG L_N=L_N_TG
x2 VDD di_spdt_ctrl_n VSS v_b v_c di_spdt_ctrl transmission_gate_lv_wo_dummy W_P=W_P_TG L_P=L_P_TG W_N=W_N_TG L_N=L_N_TG
x8 VDD di_spdt_ctrl di_spdt_ctrl_n VSS inverter_lv W_P=W_P_TG L_P=L_P_TG W_N=W_N_TG L_N=L_N_TG
.ends


* expanding   symbol:  dac_icms_cell/dac_switch.sym # of pins=6
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/dac_icms_cell/dac_switch.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/dac_icms_cell/dac_switch.sch
.subckt dac_switch VDD di_spdt_ctrl VSS v_c v_b v_a  W_P_TG=3.0u L_P_TG=0.13u W_N_TG=1.0u L_N_TG=0.13u
*.iopin v_a
*.iopin v_c
*.iopin VDD
*.iopin VSS
*.ipin di_spdt_ctrl
*.iopin v_b
x1 VDD di_spdt_ctrl VSS v_c v_a di_spdt_ctrl_n transmission_gate_lv_w_dummy W_P=W_P_TG L_P=L_P_TG W_N=W_N_TG L_N=L_N_TG W_P_D=1.0u
+ L_P_D=0.13u W_N_D=1.0u L_N_D=0.13u
x8 VDD di_spdt_ctrl di_spdt_ctrl_n VSS inverter_lv W_P=W_P_TG L_P=L_P_TG W_N=W_N_TG L_N=L_N_TG
XM1 net1 v_b VSS VSS sg13_lv_nmos w=0.5u l=0.2u ng=1 m=1
XM3 net1 v_b VDD VDD sg13_lv_pmos w=1u l=0.2u ng=1 m=1
x2 VDD di_spdt_ctrl_n VSS net1 v_c di_spdt_ctrl transmission_gate_lv_w_dummy W_P=W_P_TG L_P=L_P_TG W_N=W_N_TG L_N=L_N_TG
+ W_P_D=1.0u L_P_D=0.13u W_N_D=1.0u L_N_D=0.13u
.ends


* expanding   symbol:  transmission_gate/transmission_gate_lv_w_dummy.sym # of pins=6
** sym_path: /foss/designs/SAR_ADC_IHP/xschem/transmission_gate/transmission_gate_lv_w_dummy.sym
** sch_path: /foss/designs/SAR_ADC_IHP/xschem/transmission_gate/transmission_gate_lv_w_dummy.sch
.subckt transmission_gate_lv_w_dummy VDD di_tg_ctrl VSS v_b v_a di_tg_ctrl_n  W_P=2.0u L_P=0.13u W_N=2.0u L_N=0.13u W_P_D=1.0u
+ L_P_D=0.13u W_N_D=1.0u L_N_D=0.13u
*.iopin v_a
*.iopin v_b
*.iopin VDD
*.iopin VSS
*.ipin di_tg_ctrl
*.ipin di_tg_ctrl_n
XM1 v_a di_tg_ctrl v_b VSS sg13_lv_nmos w=W_N l=L_N ng=1 m=1
XM2 v_a di_tg_ctrl_n v_b VDD sg13_lv_pmos w=W_P l=L_P ng=1 m=1
XMdummy2 v_b di_tg_ctrl v_b VDD sg13_lv_pmos w=W_P_D l=L_P_D ng=1 m=1
XMdummy1 v_b di_tg_ctrl_n v_b VSS sg13_lv_nmos w=W_N_D l=L_N_D ng=1 m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.end
